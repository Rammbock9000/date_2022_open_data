--------------------------------------------------------------------------------
--                         ModuloCounter_56_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_56_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of ModuloCounter_56_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(5 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 55 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1718308_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1718310)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1718308_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1718308_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1718313
--                  (IntAdderAlternative_27_f250_uid1718317)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1718313 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1718313 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1718320
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1718320 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1718320 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1718323
--                   (IntAdderClassical_34_f250_uid1718325)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1718323 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1718323 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1718308
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1718308 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1718308 is
   component FPAdd_8_23_uid1718308_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1718313 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1718320 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1718323 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1718308_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1718313  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1718320  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1718323  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid1718308 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid1718308  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_56_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_56_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_56_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1718639
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1718639 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1718639 is
signal XX_m1718640 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m1718640 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m1718640 <= X ;
   YY_m1718640 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid1718643
--                   (IntAdderClassical_33_f500_uid1718645)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid1718643 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid1718643 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1718639 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid1718643 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1718639  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid1718643  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_53_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_53_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_53_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_51_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_51_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_51_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_49_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_49_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_49_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1718902_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1718904)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1718902_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1718902_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1718907
--                  (IntAdderAlternative_27_f250_uid1718911)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1718907 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1718907 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1718914
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1718914 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1718914 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1718917
--                   (IntAdderClassical_34_f250_uid1718919)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1718917 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1718917 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1718902
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1718902 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1718902 is
   component FPAdd_8_23_uid1718902_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1718907 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1718914 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1718917 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1718902_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1718907  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1718914  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1718917  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid1718902 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid1718902  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_44_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_44_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_44_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_41_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_41_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_41_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "001" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "010" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "011" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "100" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "001" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "010" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "011" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "100" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "010" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "011" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "100" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "001" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "011" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "100" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "001" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "010" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "011" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "100" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "001" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "010" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "011" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "100" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "001" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "010" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "001" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "010" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "011" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "100" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "001" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "010" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "011" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "100" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "001" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "010" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "011" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "100" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "001" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "010" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "011" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "100" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "010" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "011" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "100" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "001" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "001" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "010" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "011" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "100" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "011" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "100" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "001" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "010" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "011" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "100" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "001" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "010" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "001" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "010" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "011" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "100" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "001" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "010" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "011" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "100" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "001" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "010" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "011" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "100" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "001" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "010" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "011" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "100" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "010" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "011" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "100" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "001" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "010" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "011" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "100" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "001" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "011" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "100" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "001" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "010" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "011" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "100" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "001" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "010" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "001" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "010" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "011" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "100" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "001" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "010" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "011" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "100" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "001" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "010" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "011" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "100" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "001" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "010" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "011" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "100" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "001" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "010" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "011" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "100" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "001" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "010" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "011" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "100" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "011" when "000011",
      "000" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "100" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "001" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "010" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "000" when "000100",
      "011" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "100" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "001" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "010" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "001" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "010" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "011" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "100" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "001" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "010" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "000" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "011" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "100" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "000" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "110010" when "000000",
      "110011" when "000001",
      "000100" when "000010",
      "100100" when "000011",
      "101100" when "000100",
      "001101" when "000101",
      "000000" when "000110",
      "000001" when "000111",
      "000011" when "001000",
      "011010" when "001001",
      "000010" when "001010",
      "011000" when "001011",
      "011001" when "001100",
      "011110" when "001101",
      "001011" when "001110",
      "011101" when "001111",
      "100001" when "010000",
      "101000" when "010001",
      "000111" when "010010",
      "010111" when "010011",
      "011111" when "010100",
      "011100" when "010101",
      "001000" when "010110",
      "101011" when "010111",
      "001110" when "011000",
      "001100" when "011001",
      "100111" when "011010",
      "001001" when "011011",
      "001010" when "011100",
      "100000" when "011101",
      "000101" when "011110",
      "110100" when "011111",
      "011011" when "100000",
      "110001" when "100001",
      "101001" when "100010",
      "101010" when "100011",
      "100110" when "100100",
      "100101" when "100101",
      "101110" when "100110",
      "010010" when "100111",
      "000000" when "101000",
      "010110" when "101001",
      "010100" when "101010",
      "010011" when "101011",
      "000000" when "101100",
      "001111" when "101101",
      "010101" when "101110",
      "101111" when "101111",
      "010000" when "110000",
      "100011" when "110001",
      "010001" when "110010",
      "000000" when "110011",
      "000110" when "110100",
      "110000" when "110101",
      "100010" when "110110",
      "101101" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011110" when "000000",
      "010000" when "000001",
      "101110" when "000010",
      "000111" when "000011",
      "011011" when "000100",
      "110001" when "000101",
      "000000" when "000110",
      "101000" when "000111",
      "101011" when "001000",
      "000100" when "001001",
      "101001" when "001010",
      "010110" when "001011",
      "010111" when "001100",
      "011000" when "001101",
      "101100" when "001110",
      "000110" when "001111",
      "011001" when "010000",
      "001010" when "010001",
      "100111" when "010010",
      "010101" when "010011",
      "000010" when "010100",
      "000101" when "010101",
      "110010" when "010110",
      "011100" when "010111",
      "110000" when "011000",
      "101111" when "011001",
      "011010" when "011010",
      "110011" when "011011",
      "110100" when "011100",
      "100100" when "011101",
      "101010" when "011110",
      "010100" when "011111",
      "001101" when "100000",
      "001111" when "100001",
      "001011" when "100010",
      "001100" when "100011",
      "001001" when "100100",
      "001000" when "100101",
      "000011" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "100011" when "101001",
      "011101" when "101010",
      "000001" when "101011",
      "100101" when "101100",
      "100110" when "101101",
      "100001" when "101110",
      "010011" when "101111",
      "100000" when "110000",
      "010001" when "110001",
      "011111" when "110010",
      "000000" when "110011",
      "101101" when "110100",
      "010010" when "110101",
      "100010" when "110110",
      "001110" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "001100" when "000000",
      "001111" when "000001",
      "001101" when "000010",
      "010000" when "000011",
      "001010" when "000100",
      "011100" when "000101",
      "000000" when "000110",
      "010001" when "000111",
      "011010" when "001000",
      "100111" when "001001",
      "011011" when "001010",
      "101110" when "001011",
      "101011" when "001100",
      "101101" when "001101",
      "100000" when "001110",
      "011111" when "001111",
      "101000" when "010000",
      "001000" when "010001",
      "000000" when "010010",
      "010011" when "010011",
      "010111" when "010100",
      "010100" when "010101",
      "011101" when "010110",
      "000001" when "010111",
      "000110" when "011000",
      "010101" when "011001",
      "011110" when "011010",
      "011000" when "011011",
      "011001" when "011100",
      "000000" when "011101",
      "001011" when "011110",
      "110000" when "011111",
      "101111" when "100000",
      "000011" when "100001",
      "100110" when "100010",
      "001001" when "100011",
      "000111" when "100100",
      "100011" when "100101",
      "000100" when "100110",
      "000101" when "100111",
      "000000" when "101000",
      "000010" when "101001",
      "110001" when "101010",
      "010110" when "101011",
      "101010" when "101100",
      "101001" when "101101",
      "100100" when "101110",
      "100101" when "101111",
      "100010" when "110000",
      "100001" when "110001",
      "101100" when "110010",
      "000000" when "110011",
      "110010" when "110100",
      "010010" when "110101",
      "001110" when "110110",
      "000000" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "011111" when "000001",
      "000001" when "000010",
      "100100" when "000011",
      "100011" when "000100",
      "010001" when "000101",
      "000000" when "000110",
      "100101" when "000111",
      "010010" when "001000",
      "010011" when "001001",
      "100110" when "001010",
      "010000" when "001011",
      "011010" when "001100",
      "001111" when "001101",
      "001000" when "001110",
      "000111" when "001111",
      "011100" when "010000",
      "101110" when "010001",
      "000000" when "010010",
      "000011" when "010011",
      "000110" when "010100",
      "000100" when "010101",
      "011001" when "010110",
      "101010" when "010111",
      "101011" when "011000",
      "000010" when "011001",
      "011000" when "011010",
      "000101" when "011011",
      "011011" when "011100",
      "000000" when "011101",
      "110001" when "011110",
      "100010" when "011111",
      "100001" when "100000",
      "101111" when "100001",
      "011110" when "100010",
      "101101" when "100011",
      "101100" when "100100",
      "011101" when "100101",
      "110000" when "100110",
      "110010" when "100111",
      "000000" when "101000",
      "101001" when "101001",
      "010100" when "101010",
      "001101" when "101011",
      "010101" when "101100",
      "001110" when "101101",
      "001011" when "101110",
      "001100" when "101111",
      "001010" when "110000",
      "001001" when "110001",
      "010110" when "110010",
      "000000" when "110011",
      "010111" when "110100",
      "100111" when "110101",
      "100000" when "110110",
      "101000" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "110000" when "000000",
      "101111" when "000001",
      "101011" when "000010",
      "100101" when "000011",
      "101010" when "000100",
      "001100" when "000101",
      "000000" when "000110",
      "011001" when "000111",
      "100001" when "001000",
      "011011" when "001001",
      "001010" when "001010",
      "010011" when "001011",
      "001001" when "001100",
      "100000" when "001101",
      "011101" when "001110",
      "011000" when "001111",
      "100111" when "010000",
      "000101" when "010001",
      "000010" when "010010",
      "010000" when "010011",
      "011110" when "010100",
      "010111" when "010101",
      "010101" when "010110",
      "010100" when "010111",
      "011010" when "011000",
      "011100" when "011001",
      "000001" when "011010",
      "010110" when "011011",
      "010010" when "011100",
      "011111" when "011101",
      "101110" when "011110",
      "101101" when "011111",
      "101100" when "100000",
      "000111" when "100001",
      "100110" when "100010",
      "000110" when "100011",
      "000100" when "100100",
      "100100" when "100101",
      "000011" when "100110",
      "001110" when "100111",
      "000000" when "101000",
      "001101" when "101001",
      "100010" when "101010",
      "000000" when "101011",
      "001111" when "101100",
      "001000" when "101101",
      "010001" when "101110",
      "110100" when "101111",
      "001011" when "110000",
      "100011" when "110001",
      "101000" when "110010",
      "000000" when "110011",
      "110010" when "110100",
      "110001" when "110101",
      "110011" when "110110",
      "101001" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100010" when "000000",
      "100001" when "000001",
      "011111" when "000010",
      "001011" when "000011",
      "011110" when "000100",
      "100110" when "000101",
      "000000" when "000110",
      "011011" when "000111",
      "011101" when "001000",
      "011100" when "001001",
      "101010" when "001010",
      "010111" when "001011",
      "101100" when "001100",
      "101000" when "001101",
      "000101" when "001110",
      "001001" when "001111",
      "100000" when "010000",
      "110000" when "010001",
      "101110" when "010010",
      "011001" when "010011",
      "000100" when "010100",
      "001000" when "010101",
      "000111" when "010110",
      "000110" when "010111",
      "011010" when "011000",
      "000010" when "011001",
      "101101" when "011010",
      "000011" when "011011",
      "010110" when "011100",
      "100111" when "011101",
      "010001" when "011110",
      "010000" when "011111",
      "011000" when "100000",
      "110011" when "100001",
      "001100" when "100010",
      "110001" when "100011",
      "101111" when "100100",
      "001010" when "100101",
      "110010" when "100110",
      "000001" when "100111",
      "000000" when "101000",
      "101011" when "101001",
      "100101" when "101010",
      "101001" when "101011",
      "000000" when "101100",
      "110100" when "101101",
      "100011" when "101110",
      "001111" when "101111",
      "100100" when "110000",
      "010010" when "110001",
      "001110" when "110010",
      "000000" when "110011",
      "010100" when "110100",
      "010011" when "110101",
      "010101" when "110110",
      "001101" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "001110" when "000001",
      "010011" when "000010",
      "100101" when "000011",
      "001111" when "000100",
      "101111" when "000101",
      "000000" when "000110",
      "010000" when "000111",
      "001001" when "001000",
      "100110" when "001001",
      "101110" when "001010",
      "001000" when "001011",
      "101010" when "001100",
      "101011" when "001101",
      "000100" when "001110",
      "100010" when "001111",
      "100111" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "000010" when "010011",
      "000011" when "010100",
      "011010" when "010101",
      "011001" when "010110",
      "010101" when "010111",
      "010110" when "011000",
      "011101" when "011001",
      "001100" when "011010",
      "001101" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "001010" when "011110",
      "010100" when "011111",
      "100000" when "100000",
      "011011" when "100001",
      "011000" when "100010",
      "010111" when "100011",
      "011100" when "100100",
      "011111" when "100101",
      "000001" when "100110",
      "011110" when "100111",
      "000000" when "101000",
      "101000" when "101001",
      "101101" when "101010",
      "101100" when "101011",
      "101001" when "101100",
      "000111" when "101101",
      "100100" when "101110",
      "000110" when "101111",
      "000101" when "110000",
      "100011" when "110001",
      "001011" when "110010",
      "000000" when "110011",
      "110000" when "110100",
      "010010" when "110101",
      "100001" when "110110",
      "010001" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "011111" when "000000",
      "100000" when "000001",
      "011101" when "000010",
      "010000" when "000011",
      "011100" when "000100",
      "010111" when "000101",
      "000000" when "000110",
      "100001" when "000111",
      "101010" when "001000",
      "001111" when "001001",
      "010001" when "001010",
      "110000" when "001011",
      "010110" when "001100",
      "001100" when "001101",
      "101011" when "001110",
      "001000" when "001111",
      "011011" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "100100" when "010011",
      "100101" when "010100",
      "000101" when "010101",
      "000110" when "010110",
      "010011" when "010111",
      "010100" when "011000",
      "011010" when "011001",
      "100110" when "011010",
      "101000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "100011" when "011110",
      "010010" when "011111",
      "000010" when "100000",
      "000111" when "100001",
      "000100" when "100010",
      "000011" when "100011",
      "011001" when "100100",
      "000000" when "100101",
      "100111" when "100110",
      "000001" when "100111",
      "000000" when "101000",
      "001011" when "101001",
      "001110" when "101010",
      "001101" when "101011",
      "010101" when "101100",
      "101110" when "101101",
      "001010" when "101110",
      "101101" when "101111",
      "101100" when "110000",
      "001001" when "110001",
      "101111" when "110010",
      "000000" when "110011",
      "011000" when "110100",
      "100010" when "110101",
      "011110" when "110110",
      "101001" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000110" when "000000",
      "000011" when "000001",
      "001000" when "000010",
      "101010" when "000011",
      "000101" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "101001" when "000111",
      "100111" when "001000",
      "100110" when "001001",
      "101000" when "001010",
      "011110" when "001011",
      "100101" when "001100",
      "100100" when "001101",
      "011111" when "001110",
      "011011" when "001111",
      "000000" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "010000" when "010011",
      "010101" when "010100",
      "010001" when "010101",
      "000001" when "010110",
      "001001" when "010111",
      "000100" when "011000",
      "010100" when "011001",
      "010010" when "011010",
      "000000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "000000" when "011110",
      "000111" when "011111",
      "010011" when "100000",
      "001110" when "100001",
      "010110" when "100010",
      "001101" when "100011",
      "010111" when "100100",
      "001111" when "100101",
      "011000" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "100000" when "101001",
      "000010" when "101010",
      "100011" when "101011",
      "100010" when "101100",
      "100001" when "101101",
      "011100" when "101110",
      "011101" when "101111",
      "011010" when "110000",
      "011001" when "110001",
      "000000" when "110010",
      "000000" when "110011",
      "101011" when "110100",
      "001011" when "110101",
      "001100" when "110110",
      "001010" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "101011" when "000001",
      "100011" when "000010",
      "001011" when "000011",
      "100101" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "001010" when "000111",
      "001110" when "001000",
      "001101" when "001001",
      "001111" when "001010",
      "001001" when "001011",
      "100001" when "001100",
      "100000" when "001101",
      "011011" when "001110",
      "000101" when "001111",
      "000000" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "010111" when "010011",
      "010001" when "010100",
      "011000" when "010101",
      "101000" when "010110",
      "010000" when "010111",
      "100111" when "011000",
      "100110" when "011001",
      "000010" when "011010",
      "000000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "101001" when "011110",
      "010101" when "011111",
      "000001" when "100000",
      "000011" when "100001",
      "011001" when "100010",
      "000100" when "100011",
      "011010" when "100100",
      "010110" when "100101",
      "010100" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "001100" when "101001",
      "101010" when "101010",
      "100100" when "101011",
      "100010" when "101100",
      "010010" when "101101",
      "011110" when "101110",
      "011111" when "101111",
      "011101" when "110000",
      "011100" when "110001",
      "000000" when "110010",
      "000000" when "110011",
      "010011" when "110100",
      "001000" when "110101",
      "000111" when "110110",
      "000110" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "001001" when "000000",
      "101111" when "000001",
      "001000" when "000010",
      "100101" when "000011",
      "101010" when "000100",
      "011110" when "000101",
      "000000" when "000110",
      "000110" when "000111",
      "011100" when "001000",
      "011000" when "001001",
      "011101" when "001010",
      "011011" when "001011",
      "011010" when "001100",
      "001100" when "001101",
      "001111" when "001110",
      "000111" when "001111",
      "101001" when "010000",
      "101000" when "010001",
      "011001" when "010010",
      "010000" when "010011",
      "100010" when "010100",
      "000101" when "010101",
      "011111" when "010110",
      "010101" when "010111",
      "100000" when "011000",
      "010111" when "011001",
      "100001" when "011010",
      "010110" when "011011",
      "010010" when "011100",
      "001011" when "011101",
      "000001" when "011110",
      "101110" when "011111",
      "101100" when "100000",
      "101011" when "100001",
      "100110" when "100010",
      "100111" when "100011",
      "100100" when "100100",
      "100011" when "100101",
      "101101" when "100110",
      "110000" when "100111",
      "000000" when "101000",
      "010011" when "101001",
      "010100" when "101010",
      "001010" when "101011",
      "001110" when "101100",
      "110100" when "101101",
      "010001" when "101110",
      "000100" when "101111",
      "000010" when "110000",
      "110011" when "110001",
      "000000" when "110010",
      "000000" when "110011",
      "000011" when "110100",
      "110001" when "110101",
      "110010" when "110110",
      "001101" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "110010" when "000000",
      "100001" when "000001",
      "110000" when "000010",
      "000011" when "000011",
      "011001" when "000100",
      "000110" when "000101",
      "000000" when "000110",
      "101000" when "000111",
      "011000" when "001000",
      "010101" when "001001",
      "100100" when "001010",
      "100111" when "001011",
      "100110" when "001100",
      "101010" when "001101",
      "010011" when "001110",
      "101011" when "001111",
      "011100" when "010000",
      "011101" when "010001",
      "100101" when "010010",
      "010010" when "010011",
      "010001" when "010100",
      "101101" when "010101",
      "010110" when "010110",
      "000001" when "010111",
      "010111" when "011000",
      "010100" when "011001",
      "010000" when "011010",
      "000010" when "011011",
      "001001" when "011100",
      "101001" when "011101",
      "110001" when "011110",
      "100011" when "011111",
      "001100" when "100000",
      "001010" when "100001",
      "011110" when "100010",
      "011111" when "100011",
      "011011" when "100100",
      "011010" when "100101",
      "001011" when "100110",
      "001110" when "100111",
      "000000" when "101000",
      "000101" when "101001",
      "000100" when "101010",
      "101100" when "101011",
      "100000" when "101100",
      "001111" when "101101",
      "100010" when "101110",
      "110100" when "101111",
      "101111" when "110000",
      "001101" when "110001",
      "101110" when "110010",
      "000000" when "110011",
      "110011" when "110100",
      "000111" when "110101",
      "001000" when "110110",
      "000000" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "010001" when "000000",
      "101000" when "000001",
      "010100" when "000010",
      "000100" when "000011",
      "000010" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "100111" when "000111",
      "000011" when "001000",
      "100101" when "001001",
      "000000" when "001010",
      "100001" when "001011",
      "001110" when "001100",
      "100100" when "001101",
      "001011" when "001110",
      "011111" when "001111",
      "000000" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "001001" when "010011",
      "011010" when "010100",
      "010110" when "010101",
      "001000" when "010110",
      "011001" when "010111",
      "011000" when "011000",
      "010000" when "011001",
      "010010" when "011010",
      "000000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "010111" when "011110",
      "010011" when "011111",
      "011100" when "100000",
      "000111" when "100001",
      "011011" when "100010",
      "000000" when "100011",
      "001010" when "100100",
      "010101" when "100101",
      "011101" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "100010" when "101001",
      "001111" when "101010",
      "100011" when "101011",
      "000000" when "101100",
      "000101" when "101101",
      "100000" when "101110",
      "001101" when "101111",
      "001100" when "110000",
      "011110" when "110001",
      "000000" when "110010",
      "000000" when "110011",
      "000110" when "110100",
      "000001" when "110101",
      "100110" when "110110",
      "000000" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "010001" when "000000",
      "000111" when "000001",
      "010100" when "000010",
      "100111" when "000011",
      "100001" when "000100",
      "000000" when "000101",
      "000000" when "000110",
      "000110" when "000111",
      "100110" when "001000",
      "000100" when "001001",
      "000000" when "001010",
      "000010" when "001011",
      "100101" when "001100",
      "010010" when "001101",
      "100010" when "001110",
      "000001" when "001111",
      "000000" when "010000",
      "000000" when "010001",
      "000000" when "010010",
      "011011" when "010011",
      "001110" when "010100",
      "001100" when "010101",
      "011000" when "010110",
      "010111" when "010111",
      "010110" when "011000",
      "011100" when "011001",
      "001011" when "011010",
      "000000" when "011011",
      "000000" when "011100",
      "000000" when "011101",
      "010101" when "011110",
      "001010" when "011111",
      "001001" when "100000",
      "011110" when "100001",
      "001101" when "100010",
      "011010" when "100011",
      "011101" when "100100",
      "000000" when "100101",
      "001000" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "000011" when "101001",
      "100100" when "101010",
      "010011" when "101011",
      "000000" when "101100",
      "100011" when "101101",
      "010000" when "101110",
      "100000" when "101111",
      "011111" when "110000",
      "001111" when "110001",
      "000000" when "110010",
      "000000" when "110011",
      "101000" when "110100",
      "011001" when "110101",
      "000101" when "110110",
      "000000" when "110111",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_56_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(5 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_56_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_53_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_51_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_49_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_44_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_41_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount561_out : std_logic_vector(5 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product11_4_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product11_4_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product31_4_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product31_4_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product12_4_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product12_4_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product22_4_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product22_4_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No15_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No5_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No16_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No6_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No17_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No7_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No8_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No14_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No9_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No30_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No31_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No1_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No32_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No2_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No3_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay61No4_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No21_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No19_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No35_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No36_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay25No39_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount561_instance: ModuloCounter_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount561_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg36_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg36_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg210_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg210_out;
SharedReg166_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg166_out;
SharedReg188_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg188_out;
SharedReg232_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg254_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg254_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg210_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg188_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg254_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg166_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg188_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg188_out;
SharedReg210_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg210_out;
SharedReg232_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg254_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg254_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg210_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg254_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg36_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg36_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg166_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg188_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg188_out;
SharedReg210_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg210_out;
SharedReg232_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg254_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg254_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg210_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg254_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg36_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg62_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg88_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg114_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg140_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg166_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg188_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg188_out;
SharedReg210_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg210_out;
SharedReg232_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg254_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg254_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg210_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg254_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg609_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg609_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg609_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg609_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg422_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg445_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg468_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg468_out;
SharedReg491_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg514_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg514_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg468_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg491_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg514_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg609_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg422_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg445_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg468_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg468_out;
SharedReg491_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg514_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg514_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg468_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg491_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg514_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg609_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg609_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg422_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg445_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg468_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg468_out;
SharedReg491_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg514_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg514_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg468_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg491_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg514_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg609_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg609_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg609_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg609_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg422_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg445_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg468_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg468_out;
SharedReg491_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg514_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg514_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg468_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg491_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg514_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg609_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg630_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg651_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg651_out;
SharedReg672_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg693_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg693_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg651_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg693_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg180_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg180_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg284_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg284_out;
SharedReg282_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg282_out;
SharedReg281_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg281_out;
SharedReg281_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg281_out;
SharedReg538_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg538_out;
SharedReg433_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg433_out;
SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg276_out;
SharedReg279_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg279_out;
SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg53_out;
SharedReg438_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg438_out;
SharedReg183_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg183_out;
SharedReg442_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg442_out;
SharedReg628_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg628_out;
SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg276_out;
SharedReg186_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg186_out;
SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg364_out;
SharedReg170_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg170_out;
SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg422_out;
SharedReg620_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg620_out;
SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg422_out;
SharedReg429_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg429_out;
SharedReg432_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg432_out;
SharedReg48_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg48_out;
SharedReg616_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg616_out;
Delay25No15_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast <= Delay25No15_out;
SharedReg284_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg284_out;
SharedReg282_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg282_out;
SharedReg280_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg280_out;
SharedReg50_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg50_out;
SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg422_out;
SharedReg610_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg610_out;
SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg276_out;
SharedReg436_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg436_out;
SharedReg425_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg425_out;
SharedReg40_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg40_out;
SharedReg614_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg614_out;
SharedReg427_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg427_out;
SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg276_out;
SharedReg423_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg423_out;
SharedReg172_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg172_out;
SharedReg286_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg286_out;
SharedReg46_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg46_out;
SharedReg428_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg428_out;
SharedReg549_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg549_out;
SharedReg621_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg621_out;
SharedReg432_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg432_out;
SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg422_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg180_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg282_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg281_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg281_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg538_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg433_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg279_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg53_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg438_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg183_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg442_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg628_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg186_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg364_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg170_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg620_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg429_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg5_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg432_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg48_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg616_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay25No15_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg284_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg282_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg280_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg50_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg610_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg436_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg425_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg40_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg614_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg427_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg276_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg423_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg172_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg286_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg7_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg46_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg428_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg549_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg621_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg432_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg422_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg10_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg284_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg186_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg546_out;
SharedReg367_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg367_out;
SharedReg364_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg364_out;
SharedReg362_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg362_out;
SharedReg537_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg537_out;
SharedReg621_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg621_out;
SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg363_out;
SharedReg276_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg276_out;
SharedReg178_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg178_out;
SharedReg434_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg434_out;
SharedReg181_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg181_out;
Delay61No5_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast <= Delay61No5_out;
SharedReg629_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg629_out;
SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg363_out;
SharedReg187_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg187_out;
SharedReg358_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg358_out;
SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg167_out;
SharedReg613_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg613_out;
SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg422_out;
SharedReg610_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg610_out;
SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg609_out;
SharedReg423_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg423_out;
SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg167_out;
SharedReg429_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg429_out;
SharedReg592_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg592_out;
SharedReg364_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg364_out;
SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg363_out;
SharedReg591_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg591_out;
SharedReg166_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg166_out;
SharedReg437_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg437_out;
SharedReg625_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg625_out;
SharedReg589_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg589_out;
SharedReg426_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg426_out;
SharedReg439_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg439_out;
SharedReg56_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg56_out;
SharedReg627_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg627_out;
SharedReg439_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg439_out;
SharedReg361_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg361_out;
SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg609_out;
SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg167_out;
SharedReg276_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg276_out;
SharedReg58_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg58_out;
SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg422_out;
SharedReg277_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg277_out;
SharedReg442_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg442_out;
SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg422_out;
SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg609_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg367_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg364_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg362_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg537_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg621_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg276_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg178_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg434_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg181_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay61No5_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg629_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg187_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg358_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg613_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg610_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg23_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg423_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg429_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg592_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg364_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg363_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg591_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg166_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg437_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg625_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg22_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg589_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg426_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg439_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg56_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg627_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg439_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg361_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg167_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg276_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg25_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg58_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg277_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg442_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg422_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg609_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg27_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg450_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg450_out;
SharedReg586_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg586_out;
SharedReg446_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg446_out;
SharedReg194_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg596_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg596_out;
SharedReg72_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg72_out;
SharedReg451_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg451_out;
SharedReg381_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg381_out;
SharedReg642_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg642_out;
SharedReg455_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg455_out;
SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg445_out;
SharedReg202_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg202_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg13_out;
SharedReg295_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg295_out;
SharedReg293_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg293_out;
SharedReg292_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg292_out;
SharedReg292_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg292_out;
SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg551_out;
SharedReg456_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg456_out;
SharedReg287_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg287_out;
SharedReg290_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg290_out;
SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg79_out;
SharedReg461_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg461_out;
SharedReg205_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg205_out;
SharedReg465_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg465_out;
SharedReg649_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg649_out;
SharedReg276_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg276_out;
SharedReg208_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg208_out;
SharedReg376_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg376_out;
SharedReg192_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg192_out;
SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg445_out;
SharedReg641_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg641_out;
SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg445_out;
SharedReg452_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg452_out;
SharedReg455_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg455_out;
SharedReg74_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg74_out;
SharedReg637_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg637_out;
Delay25No16_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast <= Delay25No16_out;
SharedReg593_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg593_out;
SharedReg591_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg591_out;
SharedReg589_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg589_out;
SharedReg76_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg76_out;
SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg445_out;
SharedReg631_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg631_out;
SharedReg586_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg586_out;
SharedReg459_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg459_out;
SharedReg448_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg448_out;
SharedReg66_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg66_out;
SharedReg635_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg635_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg450_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg586_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg202_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg5_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg4_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg7_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg10_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg9_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg13_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg446_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg295_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg293_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg292_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg292_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg456_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg287_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg290_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg79_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg461_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg194_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg205_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg465_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg649_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg276_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg208_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg376_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg192_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg641_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg596_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg452_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg455_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg74_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg637_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => Delay25No16_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg593_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg591_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg589_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg76_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg445_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg72_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg631_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg586_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg459_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg448_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg66_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg635_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg451_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg381_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg642_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg455_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg462_out;
SharedReg540_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg540_out;
SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg630_out;
SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg189_out;
SharedReg287_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg287_out;
SharedReg84_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg84_out;
SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg445_out;
SharedReg288_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg288_out;
SharedReg465_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg465_out;
SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg630_out;
SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg208_out;
SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg31_out;
SharedReg558_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg558_out;
SharedReg380_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg380_out;
SharedReg376_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg376_out;
SharedReg374_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg374_out;
SharedReg550_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg550_out;
SharedReg642_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg642_out;
SharedReg375_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg375_out;
SharedReg287_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg287_out;
SharedReg200_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg200_out;
SharedReg457_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg457_out;
SharedReg203_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg203_out;
Delay61No6_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast <= Delay61No6_out;
SharedReg650_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg650_out;
SharedReg375_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg375_out;
SharedReg209_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg209_out;
SharedReg370_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg370_out;
SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg189_out;
SharedReg634_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg634_out;
SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg445_out;
SharedReg631_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg631_out;
SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg630_out;
SharedReg446_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg446_out;
SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg189_out;
SharedReg452_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg452_out;
SharedReg556_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg556_out;
SharedReg293_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg293_out;
SharedReg292_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg292_out;
SharedReg555_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg555_out;
SharedReg188_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg188_out;
SharedReg460_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg460_out;
SharedReg646_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg646_out;
SharedReg553_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg553_out;
SharedReg449_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg449_out;
SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg462_out;
SharedReg82_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg82_out;
SharedReg648_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg648_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg540_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg18_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg20_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg23_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg22_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg25_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg27_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg31_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg558_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg380_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg376_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg374_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg550_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg642_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg375_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg287_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg200_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg457_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg203_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => Delay61No6_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg650_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg375_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg209_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg370_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg634_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg631_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg287_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg630_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg446_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg189_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg452_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg556_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg293_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg292_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg555_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg188_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg460_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg84_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg646_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg553_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg449_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg462_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg82_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg648_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg288_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg465_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg557_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg557_out;
SharedReg555_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg555_out;
SharedReg291_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg291_out;
SharedReg102_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg102_out;
SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg468_out;
SharedReg652_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg652_out;
SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg322_out;
SharedReg482_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg482_out;
SharedReg471_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg471_out;
SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg92_out;
SharedReg656_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg656_out;
SharedReg473_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg473_out;
SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg322_out;
SharedReg469_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg469_out;
SharedReg216_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg216_out;
SharedReg560_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg560_out;
SharedReg98_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg98_out;
SharedReg474_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg474_out;
SharedReg309_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg309_out;
SharedReg663_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg663_out;
SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg478_out;
SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg468_out;
SharedReg224_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg224_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg13_out;
SharedReg306_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg306_out;
SharedReg304_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg304_out;
SharedReg303_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg303_out;
SharedReg303_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg303_out;
SharedReg334_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg334_out;
SharedReg479_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg479_out;
SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg322_out;
SharedReg301_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg301_out;
SharedReg105_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg105_out;
SharedReg484_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg484_out;
SharedReg227_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg227_out;
SharedReg488_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg488_out;
SharedReg670_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg670_out;
SharedReg586_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg586_out;
SharedReg230_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg230_out;
SharedReg304_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg304_out;
SharedReg214_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg214_out;
SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg468_out;
SharedReg662_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg662_out;
SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg468_out;
SharedReg475_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg475_out;
SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg478_out;
SharedReg100_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg100_out;
SharedReg658_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg658_out;
Delay25No17_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast <= Delay25No17_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg557_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg555_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg656_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg473_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg469_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg216_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg560_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg98_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg474_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg309_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg663_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg291_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg224_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg2_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg5_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg4_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg7_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg10_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg9_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg102_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg13_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg306_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg304_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg303_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg303_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg334_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg479_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg301_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg105_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg484_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg227_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg488_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg670_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg586_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg230_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg304_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg214_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg662_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg652_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg468_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg475_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg478_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg100_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg658_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => Delay25No17_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg322_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg482_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg471_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg92_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg327_out;
SharedReg326_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg326_out;
SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg210_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg210_out;
SharedReg483_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg483_out;
SharedReg667_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg667_out;
SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg387_out;
SharedReg472_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg472_out;
SharedReg485_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg485_out;
SharedReg108_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg108_out;
SharedReg669_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg669_out;
SharedReg485_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg485_out;
SharedReg552_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg552_out;
SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg651_out;
SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg211_out;
SharedReg298_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg298_out;
SharedReg110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg110_out;
SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg468_out;
SharedReg299_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg299_out;
SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg488_out;
SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg468_out;
SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg651_out;
SharedReg230_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg230_out;
SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg31_out;
SharedReg341_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg341_out;
SharedReg392_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg392_out;
SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg389_out;
SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg387_out;
SharedReg333_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg333_out;
SharedReg663_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg663_out;
SharedReg388_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg388_out;
SharedReg322_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg322_out;
SharedReg222_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg222_out;
SharedReg480_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg480_out;
SharedReg225_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg225_out;
Delay61No7_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast <= Delay61No7_out;
SharedReg671_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg671_out;
SharedReg303_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg303_out;
SharedReg231_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg231_out;
SharedReg298_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg298_out;
SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg211_out;
SharedReg655_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg655_out;
SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg468_out;
SharedReg652_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg652_out;
SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg651_out;
SharedReg469_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg469_out;
SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg211_out;
SharedReg475_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg475_out;
SharedReg390_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg390_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg327_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg669_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg485_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg552_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg298_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg110_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg299_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg488_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg230_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg18_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg20_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg23_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg22_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg25_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg27_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg210_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg31_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg341_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg392_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg389_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg333_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg663_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg388_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg322_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg222_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg483_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg480_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg225_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => Delay61No7_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg671_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg303_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg231_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg298_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg655_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg468_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg667_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg652_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg651_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg469_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg211_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg475_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg390_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg387_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg472_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg485_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg108_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg252_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg316_out;
SharedReg236_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg683_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg683_out;
SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg491_out;
SharedReg498_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg498_out;
SharedReg501_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg501_out;
SharedReg126_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg126_out;
SharedReg679_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg679_out;
SharedReg321_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg321_out;
SharedReg391_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg391_out;
SharedReg338_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg338_out;
SharedReg302_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg302_out;
SharedReg128_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg128_out;
SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg491_out;
SharedReg673_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg673_out;
SharedReg310_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg310_out;
SharedReg505_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg505_out;
SharedReg494_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg494_out;
SharedReg118_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg118_out;
SharedReg677_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg677_out;
SharedReg496_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg496_out;
SharedReg310_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg310_out;
SharedReg492_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg492_out;
SharedReg238_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg238_out;
SharedReg344_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg344_out;
SharedReg124_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg124_out;
SharedReg497_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg497_out;
SharedReg407_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg407_out;
SharedReg684_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg684_out;
SharedReg501_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg501_out;
SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg491_out;
SharedReg246_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg246_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg13_out;
SharedReg404_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg404_out;
SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg316_out;
SharedReg315_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg315_out;
SharedReg315_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg315_out;
SharedReg575_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg575_out;
SharedReg502_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg502_out;
SharedReg333_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg333_out;
SharedReg313_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg313_out;
SharedReg131_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg131_out;
SharedReg507_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg507_out;
SharedReg249_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg249_out;
SharedReg511_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg511_out;
SharedReg691_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg691_out;
SharedReg586_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg586_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg321_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg391_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg338_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg302_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg128_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg673_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg310_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg505_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg494_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg236_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg118_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg677_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg496_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg310_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg492_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg238_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg344_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg124_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg497_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg407_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg684_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg501_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg246_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg2_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg5_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg4_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg7_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg10_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg683_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg9_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg13_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg404_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg315_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg315_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg575_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg502_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg333_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg313_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg491_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg131_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg507_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg249_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg511_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg691_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg586_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg498_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg501_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg126_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg679_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg253_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg253_out;
SharedReg310_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg310_out;
SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg233_out;
SharedReg676_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg676_out;
SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg491_out;
SharedReg673_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg673_out;
SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg672_out;
SharedReg492_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg492_out;
SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg233_out;
SharedReg498_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg498_out;
SharedReg403_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg403_out;
SharedReg316_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg316_out;
SharedReg315_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg315_out;
SharedReg580_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg580_out;
SharedReg232_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg232_out;
SharedReg506_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg506_out;
SharedReg688_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg688_out;
SharedReg578_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg578_out;
SharedReg495_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg495_out;
SharedReg508_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg508_out;
SharedReg134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg134_out;
SharedReg690_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg690_out;
SharedReg508_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg508_out;
SharedReg335_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg335_out;
SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg672_out;
SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg233_out;
SharedReg396_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg396_out;
SharedReg136_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg136_out;
SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg491_out;
SharedReg397_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg397_out;
SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg511_out;
SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg491_out;
SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg672_out;
SharedReg252_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg252_out;
SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg31_out;
SharedReg341_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg341_out;
SharedReg392_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg392_out;
SharedReg402_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg402_out;
SharedReg400_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg400_out;
SharedReg574_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg574_out;
SharedReg684_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg684_out;
SharedReg401_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg401_out;
SharedReg333_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg333_out;
SharedReg244_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg244_out;
SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg503_out;
SharedReg247_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg247_out;
Delay61No8_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast <= Delay61No8_out;
SharedReg692_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg692_out;
SharedReg315_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg315_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg253_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg403_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg316_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg315_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg580_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg232_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg506_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg688_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg578_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg495_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg508_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg134_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg690_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg508_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg335_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg396_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg136_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg397_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg676_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg252_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg18_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg20_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg23_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg22_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg25_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg491_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg27_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg31_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg341_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg392_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg402_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg400_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg574_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg684_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg401_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg333_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg673_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg244_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg503_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg247_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => Delay61No8_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg692_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg315_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg672_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg492_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg233_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg498_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg350_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg350_out;
SharedReg350_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg564_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg564_out;
SharedReg525_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg525_out;
SharedReg345_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg345_out;
SharedReg348_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg348_out;
SharedReg157_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg157_out;
SharedReg530_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg530_out;
SharedReg271_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg271_out;
SharedReg534_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg534_out;
SharedReg712_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg712_out;
SharedReg345_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg345_out;
SharedReg274_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg274_out;
SharedReg415_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg415_out;
SharedReg258_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg258_out;
SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg514_out;
SharedReg704_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg704_out;
SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg514_out;
SharedReg521_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg521_out;
SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg524_out;
SharedReg152_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg152_out;
SharedReg700_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg700_out;
SharedReg409_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg409_out;
SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg353_out;
SharedReg351_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg351_out;
SharedReg314_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg314_out;
SharedReg154_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg154_out;
SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg514_out;
SharedReg694_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg694_out;
SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg410_out;
SharedReg528_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg528_out;
SharedReg517_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg517_out;
SharedReg144_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg144_out;
SharedReg698_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg698_out;
SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg519_out;
SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg410_out;
SharedReg515_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg515_out;
SharedReg260_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg260_out;
SharedReg356_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg356_out;
SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg150_out;
SharedReg520_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg520_out;
Delay19No14_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast <= Delay19No14_out;
SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg705_out;
SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg524_out;
SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg514_out;
SharedReg268_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg268_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg2_out;
SharedReg5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg5_out;
SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg9_out;
SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg13_out;
SharedReg417_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg417_out;
SharedReg351_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg351_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg350_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg712_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg345_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg274_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg415_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg258_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg704_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg521_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg564_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg152_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg700_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg409_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg353_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg351_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg314_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg154_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg694_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg525_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg528_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg517_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg144_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg698_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg519_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg410_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg515_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg260_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg356_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg150_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg345_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg520_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => Delay19No14_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg705_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg524_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg514_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg268_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg2_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg5_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg4_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg348_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg7_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg10_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg9_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg13_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg417_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg351_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg157_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg530_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg271_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg534_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg415_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg415_out;
SharedReg413_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg413_out;
SharedReg563_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg563_out;
SharedReg705_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg705_out;
SharedReg303_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg303_out;
SharedReg345_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg345_out;
SharedReg266_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg266_out;
SharedReg526_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg526_out;
SharedReg269_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg269_out;
Delay61No9_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= Delay61No9_out;
SharedReg713_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg713_out;
SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg414_out;
SharedReg275_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg275_out;
SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg410_out;
SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg255_out;
SharedReg697_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg697_out;
SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg514_out;
SharedReg694_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg694_out;
SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg693_out;
SharedReg515_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg515_out;
SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg255_out;
SharedReg521_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg521_out;
SharedReg605_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg605_out;
SharedReg415_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg415_out;
SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg414_out;
SharedReg604_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg604_out;
SharedReg254_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg254_out;
SharedReg529_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg529_out;
SharedReg709_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg709_out;
SharedReg602_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg602_out;
SharedReg518_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg518_out;
SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg531_out;
SharedReg160_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg160_out;
SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg711_out;
SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg531_out;
SharedReg577_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg577_out;
SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg693_out;
SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg255_out;
SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg410_out;
SharedReg162_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg162_out;
SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg514_out;
SharedReg411_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg411_out;
SharedReg534_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg534_out;
SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg514_out;
SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg693_out;
SharedReg274_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg274_out;
SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg23_out;
SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg27_out;
SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg31_out;
SharedReg607_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg607_out;
SharedReg572_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg572_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg415_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg413_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg713_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg275_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg697_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg694_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg515_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg563_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg521_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg605_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg415_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg414_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg604_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg254_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg529_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg709_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg602_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg705_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg518_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg160_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg711_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg531_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg577_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg255_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg410_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg162_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg303_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg411_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg534_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg514_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg693_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg274_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg18_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg20_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg23_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg22_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg345_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg25_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg27_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg31_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg607_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg572_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg266_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg526_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg269_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay61No9_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg278_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg278_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg365_out;
SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg543_out;
SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg358_out;
SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg543_out;
SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg543_out;
SharedReg48_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg48_out;
SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg537_out;
SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg586_out;
SharedReg281_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg281_out;
SharedReg625_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg625_out;
SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg358_out;
SharedReg60_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg60_out;
SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg537_out;
SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg586_out;
SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg276_out;
SharedReg538_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg538_out;
SharedReg595_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg595_out;
SharedReg166_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg166_out;
SharedReg177_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg177_out;
SharedReg166_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg166_out;
SharedReg175_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg175_out;
SharedReg46_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg46_out;
SharedReg432_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg432_out;
SharedReg369_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg369_out;
Delay25No30_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast <= Delay25No30_out;
SharedReg544_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg544_out;
SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg543_out;
SharedReg541_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg541_out;
SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg276_out;
SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg36_out;
SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg276_out;
SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg358_out;
SharedReg169_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg169_out;
SharedReg283_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg283_out;
SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg537_out;
SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg276_out;
SharedReg172_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg172_out;
SharedReg542_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg542_out;
SharedReg427_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg427_out;
SharedReg39_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg39_out;
SharedReg366_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg366_out;
SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg358_out;
SharedReg172_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg172_out;
SharedReg359_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg359_out;
SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg543_out;
SharedReg176_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg176_out;
SharedReg37_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg37_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg278_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg48_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg281_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg625_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg60_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg586_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg538_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg595_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg166_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg177_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg166_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg175_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg17_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg46_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg432_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg369_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay25No30_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg544_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg541_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg36_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg15_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg169_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg283_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg537_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg276_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg172_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg542_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg427_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg39_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg366_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg11_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg358_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg172_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg359_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg543_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg176_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg37_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg12_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg365_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No42_out);

SharedReg280_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg280_out;
SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg544_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg544_out;
SharedReg365_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg365_out;
SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg537_out;
SharedReg592_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg592_out;
SharedReg590_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg590_out;
SharedReg179_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg179_out;
SharedReg277_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg277_out;
SharedReg543_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg543_out;
SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg586_out;
SharedReg623_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg623_out;
SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg537_out;
Delay61No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast <= Delay61No_out;
SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg586_out;
SharedReg541_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg541_out;
SharedReg540_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg540_out;
SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg586_out;
SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg586_out;
SharedReg170_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg170_out;
SharedReg36_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg36_out;
SharedReg167_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg167_out;
SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg166_out;
SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg37_out;
SharedReg423_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg423_out;
SharedReg365_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg365_out;
SharedReg364_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg364_out;
SharedReg591_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg591_out;
SharedReg589_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg589_out;
SharedReg363_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg363_out;
SharedReg359_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg359_out;
SharedReg54_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg54_out;
SharedReg359_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg359_out;
SharedReg539_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg539_out;
SharedReg183_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg183_out;
SharedReg358_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg358_out;
SharedReg593_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg593_out;
SharedReg358_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg358_out;
SharedReg185_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg185_out;
SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg537_out;
SharedReg422_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg422_out;
SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg166_out;
SharedReg360_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg360_out;
SharedReg360_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg360_out;
SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg166_out;
SharedReg540_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg540_out;
SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg537_out;
SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg166_out;
SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg166_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg280_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg365_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg592_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg590_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg179_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg277_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg543_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg623_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => Delay61No_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg541_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg540_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg586_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg170_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg36_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg167_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg35_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg37_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg423_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg365_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg364_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg591_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg589_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg363_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg359_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg54_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg359_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg33_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg539_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg183_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg358_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg593_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg358_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg185_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg422_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg360_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg29_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg360_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg540_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg537_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg166_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg30_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg34_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg544_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg194_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg194_out;
SharedReg375_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg375_out;
SharedReg450_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg450_out;
SharedReg65_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg65_out;
SharedReg295_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg295_out;
SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg370_out;
SharedReg194_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg194_out;
SharedReg371_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg371_out;
SharedReg376_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg376_out;
SharedReg198_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg198_out;
SharedReg63_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg63_out;
SharedReg289_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg289_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg8_out;
SharedReg377_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg377_out;
SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg555_out;
SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg370_out;
SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg555_out;
SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg555_out;
SharedReg74_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg74_out;
SharedReg550_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg550_out;
SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg322_out;
SharedReg292_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg292_out;
SharedReg646_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg646_out;
SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg370_out;
SharedReg86_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg86_out;
SharedReg550_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg550_out;
SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg586_out;
SharedReg287_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg287_out;
SharedReg551_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg551_out;
SharedReg331_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg331_out;
SharedReg188_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg188_out;
SharedReg199_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg199_out;
SharedReg188_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg188_out;
SharedReg197_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg197_out;
SharedReg72_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg72_out;
SharedReg455_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg455_out;
SharedReg382_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg382_out;
Delay25No31_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast <= Delay25No31_out;
SharedReg377_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg377_out;
SharedReg376_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg376_out;
SharedReg374_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg374_out;
SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg586_out;
SharedReg62_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg62_out;
SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg586_out;
SharedReg287_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg287_out;
SharedReg191_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg191_out;
SharedReg592_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg592_out;
SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg586_out;
SharedReg276_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg276_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg194_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg375_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg63_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg289_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg3_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg17_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg15_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg11_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg12_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg16_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg8_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg450_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg377_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg74_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg550_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg322_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg292_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg646_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg65_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg86_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg550_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg287_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg551_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg331_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg188_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg199_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg188_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg295_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg197_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg72_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg455_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg382_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => Delay25No31_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg377_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg376_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg374_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg62_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg370_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg287_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg191_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg592_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg586_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg276_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg194_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg371_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg376_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg198_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No44_out);

SharedReg207_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg370_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg370_out;
SharedReg445_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg445_out;
SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg188_out;
SharedReg289_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg289_out;
SharedReg289_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg289_out;
SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg188_out;
SharedReg552_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg552_out;
SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg550_out;
SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg188_out;
SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg188_out;
SharedReg291_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg291_out;
SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg26_out;
SharedReg556_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg556_out;
SharedReg377_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg377_out;
SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg550_out;
SharedReg328_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg328_out;
SharedReg326_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg326_out;
SharedReg201_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg201_out;
SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg288_out;
SharedReg555_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg555_out;
SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg322_out;
SharedReg644_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg644_out;
SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg550_out;
Delay61No1_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast <= Delay61No1_out;
SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg322_out;
SharedReg553_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg553_out;
SharedReg552_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg552_out;
SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg322_out;
SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg322_out;
SharedReg192_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg192_out;
SharedReg62_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg62_out;
SharedReg189_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg189_out;
SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg188_out;
SharedReg63_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg63_out;
SharedReg446_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg446_out;
SharedReg377_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg377_out;
SharedReg293_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg293_out;
SharedReg555_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg555_out;
SharedReg553_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg553_out;
SharedReg292_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg292_out;
SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg288_out;
SharedReg80_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg80_out;
SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg288_out;
SharedReg372_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg372_out;
SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg205_out;
SharedReg287_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg287_out;
SharedReg557_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg557_out;
SharedReg358_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg358_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg370_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg291_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg35_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg33_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg29_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg30_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg34_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg26_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg445_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg556_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg377_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg328_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg326_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg201_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg555_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg644_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => Delay61No1_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg553_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg552_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg322_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg192_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg62_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg189_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg289_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg63_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg446_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg377_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg293_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg555_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg553_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg292_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg80_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg289_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg288_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg372_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg287_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg557_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg358_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg552_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg550_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg188_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg305_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg305_out;
SharedReg304_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg304_out;
SharedReg553_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg553_out;
SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg550_out;
SharedReg88_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg88_out;
SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg322_out;
SharedReg298_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg298_out;
SharedReg213_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg213_out;
SharedReg556_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg556_out;
SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg322_out;
SharedReg287_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg287_out;
SharedReg216_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg216_out;
SharedReg388_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg388_out;
SharedReg473_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg473_out;
SharedReg91_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg91_out;
SharedReg306_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg306_out;
SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg383_out;
SharedReg216_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg216_out;
SharedReg384_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg384_out;
SharedReg389_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg389_out;
SharedReg220_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg220_out;
SharedReg89_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg89_out;
SharedReg300_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg300_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg8_out;
SharedReg390_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg390_out;
SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg338_out;
SharedReg370_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg370_out;
SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg338_out;
SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg100_out;
SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg383_out;
SharedReg333_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg333_out;
SharedReg303_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg303_out;
SharedReg667_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg667_out;
SharedReg298_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg298_out;
SharedReg112_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg112_out;
SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg383_out;
SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg550_out;
SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg322_out;
SharedReg384_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg384_out;
SharedReg319_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg319_out;
SharedReg210_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg210_out;
SharedReg221_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg221_out;
SharedReg210_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg210_out;
SharedReg219_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg219_out;
SharedReg98_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg98_out;
SharedReg478_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg478_out;
SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg395_out;
Delay25No32_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast <= Delay25No32_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg305_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg304_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg287_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg216_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg388_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg473_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg91_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg306_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg216_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg384_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg389_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg553_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg220_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg89_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg300_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg3_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg17_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg15_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg11_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg12_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg16_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg8_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg390_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg370_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg338_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg100_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg333_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg303_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg88_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg667_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg298_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg112_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg383_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg550_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg384_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg319_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg210_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg221_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg210_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg219_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg98_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg478_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg395_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => Delay25No32_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg298_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg213_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg556_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg322_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No46_out);

SharedReg389_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg389_out;
SharedReg387_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg387_out;
SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg326_out;
SharedReg323_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg323_out;
SharedReg106_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg106_out;
SharedReg299_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg299_out;
SharedReg385_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg385_out;
SharedReg227_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg227_out;
SharedReg298_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg298_out;
SharedReg391_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg391_out;
SharedReg370_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg370_out;
SharedReg229_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg229_out;
SharedReg383_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg383_out;
SharedReg468_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg468_out;
SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg210_out;
SharedReg300_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg300_out;
SharedReg300_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg300_out;
SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg210_out;
SharedReg335_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg335_out;
SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg333_out;
SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg210_out;
SharedReg302_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg302_out;
SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg26_out;
SharedReg339_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg339_out;
SharedReg390_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg390_out;
SharedReg550_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg550_out;
SharedReg317_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg317_out;
SharedReg315_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg315_out;
SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg223_out;
SharedReg299_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg299_out;
SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg338_out;
SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg333_out;
SharedReg665_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg665_out;
SharedReg383_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg383_out;
Delay61No2_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast <= Delay61No2_out;
SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg333_out;
SharedReg387_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg387_out;
SharedReg386_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg386_out;
SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg333_out;
SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg333_out;
SharedReg214_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg214_out;
SharedReg88_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg88_out;
SharedReg211_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg211_out;
SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg210_out;
SharedReg89_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg89_out;
SharedReg469_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg469_out;
SharedReg305_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg305_out;
SharedReg327_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg327_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg389_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg387_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg370_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg229_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg383_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg468_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg300_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg300_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg335_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg326_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg302_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg19_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg21_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg35_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg33_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg29_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg30_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg34_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg323_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg26_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg339_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg390_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg550_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg317_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg315_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg223_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg299_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg338_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg106_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg665_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg383_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => Delay61No2_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg387_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg386_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg333_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg214_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg88_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg299_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg211_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg210_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg89_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg469_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg305_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg327_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg385_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg227_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg298_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg391_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg333_out;
SharedReg397_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg355_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg355_out;
SharedReg232_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg243_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg243_out;
SharedReg232_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg232_out;
SharedReg241_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg241_out;
SharedReg124_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg124_out;
SharedReg501_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg501_out;
SharedReg408_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg408_out;
SharedReg585_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg585_out;
SharedReg403_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg403_out;
SharedReg402_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg402_out;
SharedReg336_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg336_out;
SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg333_out;
SharedReg114_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg114_out;
SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg310_out;
SharedReg396_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg396_out;
SharedReg235_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg235_out;
SharedReg339_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg339_out;
SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg310_out;
SharedReg298_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg298_out;
SharedReg238_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg238_out;
SharedReg579_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg579_out;
SharedReg496_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg496_out;
SharedReg117_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg117_out;
SharedReg404_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg404_out;
SharedReg574_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg574_out;
SharedReg238_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg238_out;
SharedReg575_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg575_out;
SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg580_out;
SharedReg242_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg242_out;
SharedReg115_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg115_out;
SharedReg398_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg398_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg8_out;
SharedReg581_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg581_out;
SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg580_out;
SharedReg298_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg298_out;
SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg580_out;
SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg580_out;
SharedReg126_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg126_out;
SharedReg396_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg396_out;
SharedReg574_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg574_out;
SharedReg315_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg315_out;
SharedReg688_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg688_out;
SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg310_out;
SharedReg138_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg138_out;
SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg333_out;
SharedReg550_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg550_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg585_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg403_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg402_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg336_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg114_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg396_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg235_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg339_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg355_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg298_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg238_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg579_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg496_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg117_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg404_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg574_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg238_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg575_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg232_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg242_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg115_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg398_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg3_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg17_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg15_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg11_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg12_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg243_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg16_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg8_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg581_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg298_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg580_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg126_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg396_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg574_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg232_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg315_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg688_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg310_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg138_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg333_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg550_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg241_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg124_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg501_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg408_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No48_out);

SharedReg399_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg399_out;
SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg574_out;
SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg574_out;
SharedReg236_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg114_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg233_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg233_out;
SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg232_out;
SharedReg115_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg115_out;
SharedReg492_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg492_out;
SharedReg317_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg317_out;
SharedReg316_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg316_out;
SharedReg580_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg580_out;
SharedReg578_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg578_out;
SharedReg315_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg315_out;
SharedReg311_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg311_out;
SharedReg132_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg132_out;
SharedReg397_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg397_out;
SharedReg576_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg576_out;
SharedReg249_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg249_out;
SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg396_out;
SharedReg582_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg582_out;
SharedReg383_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg383_out;
SharedReg251_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg251_out;
SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg574_out;
SharedReg491_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg491_out;
SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg232_out;
SharedReg398_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg398_out;
SharedReg398_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg398_out;
SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg232_out;
SharedReg348_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg348_out;
SharedReg345_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg345_out;
SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg232_out;
SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg232_out;
SharedReg400_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg400_out;
SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg26_out;
SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg352_out;
SharedReg581_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg581_out;
SharedReg383_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg383_out;
SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg352_out;
SharedReg350_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg350_out;
SharedReg245_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg245_out;
SharedReg311_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg311_out;
SharedReg580_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg580_out;
SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg574_out;
SharedReg686_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg686_out;
SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg396_out;
Delay61No3_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast <= Delay61No3_out;
SharedReg310_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg310_out;
SharedReg400_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg400_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg399_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg316_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg580_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg578_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg315_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg311_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg132_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg397_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg576_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg249_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg582_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg383_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg251_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg491_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg398_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg398_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg348_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg236_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg345_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg400_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg19_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg21_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg35_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg33_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg29_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg30_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg114_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg34_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg26_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg581_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg383_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg350_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg245_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg311_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg580_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg233_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg574_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg686_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg396_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => Delay61No3_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg310_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg400_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg232_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg115_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg492_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg317_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg410_out;
SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg569_out;
SharedReg152_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg152_out;
SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg598_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg598_out;
SharedReg350_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg350_out;
SharedReg709_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg709_out;
SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg410_out;
SharedReg164_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg164_out;
SharedReg383_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg383_out;
SharedReg598_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg598_out;
SharedReg345_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg345_out;
SharedReg564_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg564_out;
SharedReg608_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg608_out;
SharedReg254_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg254_out;
SharedReg265_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg265_out;
SharedReg254_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg254_out;
SharedReg263_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg263_out;
SharedReg150_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg150_out;
SharedReg524_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg524_out;
SharedReg421_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg421_out;
SharedReg357_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg357_out;
SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg570_out;
SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg569_out;
SharedReg578_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg578_out;
SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg410_out;
SharedReg140_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg140_out;
SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg410_out;
SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg563_out;
SharedReg257_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg257_out;
SharedReg352_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg352_out;
SharedReg345_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg345_out;
SharedReg310_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg310_out;
SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg260_out;
SharedReg603_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg603_out;
SharedReg519_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg519_out;
SharedReg143_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg143_out;
SharedReg571_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg571_out;
SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg563_out;
SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg260_out;
SharedReg564_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg564_out;
SharedReg604_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg604_out;
SharedReg264_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg264_out;
SharedReg141_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg141_out;
SharedReg412_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg412_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg17_out;
SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg15_out;
SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg16_out;
SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg8_out;
SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg570_out;
SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg569_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg383_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg598_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg345_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg564_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg608_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg254_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg265_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg254_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg263_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg150_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg524_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg421_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg357_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg578_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg140_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg152_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg257_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg352_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg345_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg310_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg603_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg519_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg143_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg571_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg563_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg260_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg564_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg604_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg264_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg141_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg412_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg3_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg17_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg15_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg598_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg11_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg12_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg16_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg8_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg569_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg350_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg709_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg410_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg164_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No50_out);

SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg563_out;
SharedReg605_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg605_out;
SharedReg603_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg603_out;
SharedReg267_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg267_out;
SharedReg575_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg575_out;
SharedReg389_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg389_out;
SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg598_out;
SharedReg707_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg707_out;
SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg563_out;
Delay61No4_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= Delay61No4_out;
SharedReg333_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg333_out;
SharedReg567_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg348_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg348_out;
SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg598_out;
SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg563_out;
SharedReg258_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg258_out;
SharedReg140_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg140_out;
SharedReg255_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg255_out;
SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg254_out;
SharedReg141_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg141_out;
SharedReg515_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg515_out;
SharedReg352_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg352_out;
SharedReg415_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg415_out;
SharedReg604_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg604_out;
SharedReg413_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg413_out;
SharedReg579_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg579_out;
SharedReg411_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg411_out;
SharedReg158_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg158_out;
SharedReg564_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg564_out;
SharedReg600_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg600_out;
SharedReg271_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg271_out;
SharedReg345_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg345_out;
SharedReg606_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg606_out;
SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg396_out;
SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg273_out;
SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg598_out;
SharedReg514_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg514_out;
SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg254_out;
SharedReg565_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg565_out;
SharedReg565_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg565_out;
SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg254_out;
SharedReg601_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg601_out;
SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg598_out;
SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg254_out;
SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg254_out;
SharedReg413_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg413_out;
SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg35_out;
SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg33_out;
SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg34_out;
SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg26_out;
SharedReg605_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg605_out;
SharedReg416_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg416_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg605_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg333_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg348_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg258_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg140_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg255_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg141_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg603_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg515_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg352_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg415_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg604_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg413_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg579_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg411_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg158_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg564_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg600_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg267_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg271_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg345_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg606_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg396_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg514_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg565_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg565_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg575_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg601_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg254_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg413_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg19_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg21_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg35_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg33_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg389_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg29_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg30_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg34_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg26_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg605_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg416_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg598_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg707_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg563_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay61No4_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No52_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg747_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg747_out;
SharedReg748_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg748_out;
SharedReg749_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg749_out;
SharedReg750_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg750_out;
SharedReg751_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg751_out;
SharedReg752_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg752_out;
SharedReg714_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg714_out;
SharedReg862_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg862_out;
SharedReg858_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg858_out;
SharedReg804_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg804_out;
SharedReg763_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg763_out;
SharedReg718_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg718_out;
SharedReg809_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg809_out;
SharedReg720_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg720_out;
SharedReg842_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg842_out;
SharedReg816_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg816_out;
SharedReg427_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg427_out;
SharedReg426_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg426_out;
SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg843_out;
SharedReg724_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg725_out;
SharedReg847_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg847_out;
SharedReg753_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg753_out;
SharedReg754_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg758_out;
SharedReg759_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg759_out;
SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg843_out;
SharedReg727_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg727_out;
SharedReg728_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg728_out;
SharedReg729_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg729_out;
SharedReg730_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg730_out;
SharedReg731_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg731_out;
SharedReg732_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg732_out;
SharedReg808_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg808_out;
SharedReg614_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg614_out;
SharedReg734_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg734_out;
SharedReg735_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg735_out;
SharedReg736_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg736_out;
SharedReg172_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg172_out;
SharedReg738_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg738_out;
SharedReg739_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg739_out;
SharedReg740_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg740_out;
SharedReg784_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg784_out;
SharedReg741_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg741_out;
SharedReg786_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg786_out;
SharedReg787_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg787_out;
SharedReg48_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg48_out;
SharedReg743_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg743_out;
SharedReg736_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg744_out;
SharedReg745_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg745_out;
SharedReg746_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg746_out;
SharedReg822_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg822_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg747_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg748_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg763_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg718_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg809_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg720_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg842_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg816_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg427_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg426_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg724_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg749_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg725_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg847_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg753_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg754_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg755_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg756_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg757_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg758_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg759_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg843_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg750_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg727_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg728_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg729_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg730_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg731_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg732_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg808_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg614_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg734_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg735_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg751_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg736_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg172_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg738_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg739_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg740_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg784_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg741_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg786_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg787_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg48_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg752_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg743_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg736_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg744_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg745_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg746_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg822_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg714_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg862_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg858_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg804_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No52_out);

SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg168_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg166_out;
SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg37_out;
SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg167_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg36_out;
SharedReg422_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg422_out;
SharedReg609_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg609_out;
SharedReg609_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg609_out;
SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg39_out;
SharedReg171_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg171_out;
SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg425_out;
SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg42_out;
SharedReg613_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg613_out;
SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg425_out;
SharedReg829_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg829_out;
SharedReg815_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg815_out;
SharedReg616_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg616_out;
SharedReg172_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg172_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg44_out;
SharedReg617_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg617_out;
SharedReg169_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg169_out;
SharedReg435_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg435_out;
SharedReg41_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg41_out;
SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg39_out;
SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg39_out;
SharedReg615_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg615_out;
SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg40_out;
SharedReg637_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg637_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg36_out;
SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg166_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg36_out;
SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg167_out;
SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg36_out;
SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg167_out;
SharedReg613_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg613_out;
SharedReg813_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg813_out;
SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg43_out;
SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg40_out;
SharedReg428_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg428_out;
SharedReg781_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg781_out;
SharedReg173_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg173_out;
SharedReg46_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg46_out;
SharedReg174_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg174_out;
SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg44_out;
SharedReg45_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg45_out;
SharedReg619_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg619_out;
SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg38_out;
SharedReg788_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg788_out;
SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg49_out;
SharedReg451_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg451_out;
SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg166_out;
SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg166_out;
SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg38_out;
SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg425_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg171_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg42_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg613_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg829_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg815_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg616_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg172_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg168_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg617_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg169_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg435_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg41_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg39_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg615_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg637_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg613_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg813_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg43_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg40_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg37_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg428_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg781_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg173_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg46_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg174_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg44_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg45_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg619_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg788_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg167_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg49_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg451_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg166_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg38_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg425_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg36_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg422_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg609_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg609_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No54_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg784_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg784_out;
SharedReg741_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg741_out;
SharedReg786_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg786_out;
SharedReg787_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg787_out;
SharedReg74_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg74_out;
SharedReg743_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg743_out;
SharedReg736_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg744_out;
SharedReg745_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg745_out;
SharedReg746_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg746_out;
SharedReg822_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg822_out;
SharedReg747_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg747_out;
SharedReg748_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg748_out;
SharedReg749_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg749_out;
SharedReg750_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg750_out;
SharedReg751_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg751_out;
SharedReg752_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg752_out;
SharedReg714_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg714_out;
SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg862_out;
SharedReg858_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg858_out;
SharedReg804_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg804_out;
SharedReg763_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg763_out;
SharedReg718_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg718_out;
SharedReg809_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg809_out;
SharedReg720_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg720_out;
SharedReg842_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg842_out;
SharedReg816_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg816_out;
SharedReg450_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg450_out;
SharedReg449_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg449_out;
SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg862_out;
SharedReg724_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg725_out;
SharedReg847_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg847_out;
SharedReg191_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg191_out;
SharedReg798_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg798_out;
SharedReg799_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg799_out;
SharedReg65_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg65_out;
SharedReg801_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg802_out;
SharedReg66_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg66_out;
SharedReg658_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg658_out;
SharedReg62_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg62_out;
SharedReg188_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg188_out;
SharedReg774_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg774_out;
SharedReg189_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg189_out;
SharedReg776_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg776_out;
SharedReg189_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg189_out;
SharedReg808_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg808_out;
SharedReg733_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg733_out;
SharedReg778_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg778_out;
SharedReg759_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg759_out;
SharedReg679_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg679_out;
SharedReg196_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg196_out;
SharedReg851_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg851_out;
SharedReg782_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg783_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg784_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg741_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg822_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg747_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg748_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg749_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg750_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg751_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg752_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg714_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg858_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg786_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg804_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg763_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg718_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg809_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg720_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg842_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg816_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg450_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg449_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg787_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg724_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg725_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg847_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg191_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg798_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg799_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg65_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg801_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg802_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg66_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg74_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg658_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg62_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg188_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg774_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg189_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg776_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg189_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg808_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg733_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg778_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg743_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg759_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg679_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg196_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg851_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg782_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg783_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg736_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg744_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg745_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg746_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No54_out);

SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg71_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg71_out;
SharedReg640_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg640_out;
SharedReg64_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg64_out;
SharedReg788_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg788_out;
SharedReg75_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg75_out;
SharedReg474_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg474_out;
SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg188_out;
SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg188_out;
SharedReg64_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg64_out;
SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg448_out;
SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg65_out;
SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg63_out;
SharedReg190_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg190_out;
SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg188_out;
SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg63_out;
SharedReg189_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg189_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg62_out;
SharedReg445_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg445_out;
SharedReg630_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg630_out;
SharedReg630_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg630_out;
SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg65_out;
SharedReg193_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg193_out;
SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg448_out;
SharedReg68_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg68_out;
SharedReg634_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg634_out;
SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg448_out;
SharedReg829_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg829_out;
SharedReg815_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg815_out;
SharedReg468_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg468_out;
SharedReg194_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg194_out;
SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg70_out;
SharedReg638_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg638_out;
SharedReg797_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg797_out;
SharedReg458_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg458_out;
SharedReg67_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg67_out;
SharedReg800_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg800_out;
SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg65_out;
SharedReg636_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg636_out;
SharedReg803_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg803_out;
SharedReg845_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg845_out;
SharedReg772_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg772_out;
SharedReg773_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg773_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg62_out;
SharedReg775_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg775_out;
SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg62_out;
SharedReg777_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg777_out;
SharedReg631_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg631_out;
SharedReg192_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg192_out;
SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg69_out;
SharedReg92_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg92_out;
SharedReg845_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg845_out;
SharedReg781_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg781_out;
SharedReg454_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg454_out;
SharedReg72_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg72_out;
SharedReg196_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg196_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg190_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg63_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg189_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg445_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg630_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg640_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg630_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg193_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg68_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg634_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg448_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg829_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg815_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg468_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg64_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg194_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg70_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg638_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg797_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg458_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg67_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg800_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg65_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg636_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg803_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg788_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg845_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg772_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg773_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg775_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg62_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg777_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg631_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg192_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg69_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg75_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg92_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg845_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg781_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg454_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg72_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg196_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg474_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg188_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg64_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No56_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg776_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg776_out;
SharedReg211_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg808_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg808_out;
SharedReg733_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg733_out;
SharedReg778_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg778_out;
SharedReg759_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg759_out;
SharedReg814_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg814_out;
SharedReg218_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg218_out;
SharedReg851_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg851_out;
SharedReg782_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg783_out;
SharedReg784_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg784_out;
SharedReg741_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg741_out;
SharedReg786_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg786_out;
SharedReg787_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg787_out;
SharedReg100_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg100_out;
SharedReg743_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg743_out;
SharedReg736_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg744_out;
SharedReg745_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg745_out;
SharedReg746_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg746_out;
SharedReg822_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg822_out;
SharedReg747_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg747_out;
SharedReg748_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg748_out;
SharedReg749_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg749_out;
SharedReg750_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg750_out;
SharedReg751_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg751_out;
SharedReg752_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg752_out;
SharedReg714_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg714_out;
SharedReg744_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg744_out;
SharedReg858_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg858_out;
SharedReg804_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg804_out;
SharedReg763_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg763_out;
SharedReg215_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg215_out;
SharedReg654_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg654_out;
SharedReg844_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg844_out;
SharedReg721_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg721_out;
SharedReg816_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg816_out;
SharedReg722_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg722_out;
SharedReg814_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg814_out;
SharedReg862_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg862_out;
SharedReg216_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg216_out;
SharedReg770_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg770_out;
SharedReg853_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg853_out;
SharedReg753_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg753_out;
SharedReg754_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg758_out;
SharedReg495_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg495_out;
SharedReg760_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg760_out;
SharedReg727_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg727_out;
SharedReg848_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg848_out;
SharedReg806_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg806_out;
SharedReg651_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg651_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg776_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg783_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg784_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg741_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg786_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg787_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg100_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg743_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg736_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg744_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg745_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg808_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg746_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg822_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg747_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg748_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg749_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg750_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg751_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg752_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg714_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg744_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg733_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg858_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg804_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg763_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg215_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg654_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg844_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg721_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg816_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg722_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg814_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg778_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg862_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg216_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg770_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg853_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg753_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg754_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg755_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg756_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg757_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg758_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg759_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg495_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg760_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg727_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg848_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg806_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg651_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg814_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg218_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg851_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg782_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No56_out);

SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg777_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg777_out;
SharedReg652_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg652_out;
SharedReg214_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg214_out;
SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg95_out;
SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg521_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg521_out;
SharedReg781_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg781_out;
SharedReg477_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg477_out;
SharedReg98_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg98_out;
SharedReg218_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg218_out;
SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg96_out;
SharedReg97_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg97_out;
SharedReg661_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg661_out;
SharedReg90_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg90_out;
SharedReg788_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg788_out;
SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg101_out;
SharedReg497_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg497_out;
SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg210_out;
SharedReg90_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg90_out;
SharedReg471_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg471_out;
SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg91_out;
SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg89_out;
SharedReg212_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg212_out;
SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg210_out;
SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg89_out;
SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg211_out;
SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg88_out;
SharedReg232_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg232_out;
SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg651_out;
SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg651_out;
SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg91_out;
SharedReg764_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg764_out;
SharedReg809_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg809_out;
SharedReg654_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg654_out;
SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg91_out;
SharedReg472_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg472_out;
SharedReg94_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg94_out;
SharedReg475_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg475_out;
SharedReg672_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg672_out;
SharedReg769_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg769_out;
SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg96_out;
SharedReg659_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg659_out;
SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg103_out;
SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg656_out;
SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg656_out;
SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg656_out;
SharedReg213_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg213_out;
SharedReg472_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg472_out;
SharedReg815_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg815_out;
SharedReg140_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg140_out;
SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg651_out;
SharedReg468_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg468_out;
SharedReg468_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg468_out;
SharedReg855_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg855_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg777_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg218_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg97_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg661_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg90_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg788_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg101_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg497_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg652_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg90_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg471_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg212_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg210_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg89_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg211_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg88_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg232_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg214_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg764_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg809_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg654_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg91_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg472_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg94_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg475_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg95_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg672_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg769_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg96_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg659_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg103_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg656_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg213_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg472_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg118_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg815_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg140_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg651_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg468_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg468_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg855_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg521_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg781_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg477_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg98_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No58_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg237_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg237_out;
SharedReg114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg114_out;
SharedReg233_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg233_out;
SharedReg232_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg117_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg117_out;
SharedReg88_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg88_out;
SharedReg238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg238_out;
SharedReg238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg238_out;
SharedReg471_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg471_out;
SharedReg652_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg652_out;
SharedReg651_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg651_out;
SharedReg677_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg677_out;
SharedReg651_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg651_out;
SharedReg677_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg677_out;
SharedReg653_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg653_out;
SharedReg675_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg675_out;
SharedReg816_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg816_out;
SharedReg815_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg815_out;
SharedReg714_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg714_out;
SharedReg763_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg763_out;
SharedReg804_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg804_out;
SharedReg844_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg844_out;
SharedReg858_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg858_out;
SharedReg738_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg738_out;
SharedReg731_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg731_out;
SharedReg732_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg732_out;
SharedReg774_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg774_out;
SharedReg717_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg717_out;
SharedReg740_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg740_out;
SharedReg734_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg734_out;
SharedReg808_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg808_out;
SharedReg739_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg739_out;
SharedReg736_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg736_out;
SharedReg850_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg850_out;
SharedReg853_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg853_out;
SharedReg722_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg722_out;
SharedReg801_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg801_out;
SharedReg751_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg751_out;
SharedReg750_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg750_out;
SharedReg841_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg841_out;
SharedReg759_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg759_out;
SharedReg748_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg748_out;
SharedReg749_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg749_out;
SharedReg838_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg838_out;
SharedReg802_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg802_out;
SharedReg753_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg753_out;
SharedReg752_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg752_out;
SharedReg721_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg721_out;
SharedReg770_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg770_out;
SharedReg747_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg747_out;
SharedReg798_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg798_out;
SharedReg799_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg799_out;
SharedReg716_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg716_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_53_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg237_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg651_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg677_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg651_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg677_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg653_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg675_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg816_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg815_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg714_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg763_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg233_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg804_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg844_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg858_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg738_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg731_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg732_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg774_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg717_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg740_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg734_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg232_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg808_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg739_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg736_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg850_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg853_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg722_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg801_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg751_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg750_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg841_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg117_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg759_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg748_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg749_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg838_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg802_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg753_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg752_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg721_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg770_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg747_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg88_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg798_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg799_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg716_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_6 => SharedReg238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg238_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg471_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg652_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product4_3_impl_0_LUT_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No58_out);

SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg124_out;
SharedReg233_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg233_out;
SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg240_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg240_out;
SharedReg121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg121_out;
SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg117_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg115_out;
SharedReg232_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg232_out;
SharedReg144_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg144_out;
SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg115_out;
SharedReg234_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg234_out;
SharedReg89_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg89_out;
SharedReg129_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg129_out;
SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg117_out;
SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg119_out;
SharedReg120_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg120_out;
SharedReg122_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg122_out;
SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg117_out;
SharedReg210_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg210_out;
SharedReg239_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg239_out;
SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg114_out;
SharedReg233_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg233_out;
SharedReg676_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg676_out;
SharedReg680_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg680_out;
SharedReg469_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg469_out;
SharedReg678_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg678_out;
SharedReg469_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg469_out;
SharedReg672_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg672_out;
SharedReg504_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg504_out;
SharedReg498_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg498_out;
SharedReg495_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg495_out;
SharedReg675_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg675_out;
SharedReg680_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg680_out;
SharedReg672_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg672_out;
SharedReg520_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg520_out;
SharedReg764_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg764_out;
SharedReg809_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg809_out;
SharedReg781_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg781_out;
SharedReg772_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg772_out;
SharedReg775_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg775_out;
SharedReg761_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg761_out;
SharedReg773_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg773_out;
SharedReg813_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg813_out;
SharedReg769_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg769_out;
SharedReg800_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg800_out;
SharedReg840_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg840_out;
SharedReg839_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg839_out;
SharedReg803_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg803_out;
SharedReg837_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg837_out;
SharedReg796_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg796_out;
SharedReg760_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg760_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_53_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg144_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg234_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg89_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg129_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg119_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg120_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg122_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg124_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg210_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg239_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg233_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg676_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg680_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg469_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg678_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg469_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg672_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg233_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg504_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg498_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg495_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg675_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg680_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg672_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg520_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg764_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg809_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg781_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg114_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg772_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg775_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg761_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg773_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg813_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg769_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg800_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg840_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg839_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg803_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg240_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg837_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg796_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg760_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_6 => SharedReg121_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg117_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg115_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg232_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product4_3_impl_1_LUT_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No60_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg731_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg731_out;
SharedReg732_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg732_out;
SharedReg808_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg808_out;
SharedReg656_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg656_out;
SharedReg734_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg734_out;
SharedReg850_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg850_out;
SharedReg518_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg518_out;
SharedReg216_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg216_out;
SharedReg738_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg738_out;
SharedReg739_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg739_out;
SharedReg740_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg740_out;
SharedReg448_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg448_out;
SharedReg838_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg838_out;
SharedReg632_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg632_out;
SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg630_out;
SharedReg841_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg841_out;
SharedReg631_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg631_out;
SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg630_out;
SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg630_out;
SharedReg62_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg62_out;
SharedReg716_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg716_out;
SharedReg717_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg717_out;
SharedReg805_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg805_out;
SharedReg719_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg719_out;
SharedReg861_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg861_out;
SharedReg194_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg194_out;
SharedReg66_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg66_out;
SharedReg722_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg722_out;
SharedReg815_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg815_out;
SharedReg651_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg651_out;
SharedReg196_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg196_out;
SharedReg770_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg770_out;
SharedReg771_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg771_out;
SharedReg718_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg718_out;
SharedReg809_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg809_out;
SharedReg720_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg720_out;
SharedReg842_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg842_out;
SharedReg816_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg816_out;
SharedReg473_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg473_out;
SharedReg472_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg472_out;
SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg862_out;
SharedReg724_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg725_out;
SharedReg847_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg847_out;
SharedReg213_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg213_out;
SharedReg798_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg798_out;
SharedReg799_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg799_out;
SharedReg91_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg91_out;
SharedReg801_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg802_out;
SharedReg656_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg656_out;
SharedReg714_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg714_out;
SharedReg88_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg88_out;
SharedReg210_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg210_out;
SharedReg774_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg774_out;
SharedReg211_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg211_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg731_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg732_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg740_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg448_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg838_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg632_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg841_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg631_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg630_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg62_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg808_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg716_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg717_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg805_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg719_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg861_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg194_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg66_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg722_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg815_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg651_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg656_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg196_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg770_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg771_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg718_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg809_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg720_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg842_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg816_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg473_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg472_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg734_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg724_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg725_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg847_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg213_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg798_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg799_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg91_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg801_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg802_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg850_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg656_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg714_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg88_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg210_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg774_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg211_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg518_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg216_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg738_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg739_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No60_out);

SharedReg88_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg211_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg655_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg655_out;
SharedReg813_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg813_out;
SharedReg95_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg95_out;
SharedReg659_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg659_out;
SharedReg815_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg815_out;
SharedReg781_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg781_out;
SharedReg217_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg217_out;
SharedReg98_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg98_out;
SharedReg218_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg218_out;
SharedReg837_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg837_out;
SharedReg446_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg446_out;
SharedReg839_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg839_out;
SharedReg840_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg840_out;
SharedReg446_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg446_out;
SharedReg796_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg796_out;
SharedReg760_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg760_out;
SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg863_out;
SharedReg761_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg761_out;
SharedReg188_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg188_out;
SharedReg63_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg63_out;
SharedReg447_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg447_out;
SharedReg636_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg636_out;
SharedReg631_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg631_out;
SharedReg766_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg766_out;
SharedReg767_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg767_out;
SharedReg455_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg455_out;
SharedReg452_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg452_out;
SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg863_out;
SharedReg769_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg769_out;
SharedReg198_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg198_out;
SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg70_out;
SharedReg215_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg215_out;
SharedReg471_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg471_out;
SharedReg94_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg94_out;
SharedReg655_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg655_out;
SharedReg471_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg471_out;
SharedReg829_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg829_out;
SharedReg815_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg815_out;
SharedReg491_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg491_out;
SharedReg216_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg216_out;
SharedReg96_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg96_out;
SharedReg659_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg659_out;
SharedReg797_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg797_out;
SharedReg481_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg481_out;
SharedReg93_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg93_out;
SharedReg800_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg800_out;
SharedReg91_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg91_out;
SharedReg657_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg657_out;
SharedReg803_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg803_out;
SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg140_out;
SharedReg772_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg772_out;
SharedReg773_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg773_out;
SharedReg88_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg88_out;
SharedReg775_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg775_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg218_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg837_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg446_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg839_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg840_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg446_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg796_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg760_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg761_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg655_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg188_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg63_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg447_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg636_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg631_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg766_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg767_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg455_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg452_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg813_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg769_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg198_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg70_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg215_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg471_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg94_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg655_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg471_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg829_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg815_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg95_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg491_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg216_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg96_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg659_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg797_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg481_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg93_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg800_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg91_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg657_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg659_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg803_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg140_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg772_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg773_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg88_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg775_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg815_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg781_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg217_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg98_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product11_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_3_impl_out,
                 X => Delay1No62_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg754_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg758_out;
SharedReg759_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg759_out;
SharedReg815_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg815_out;
SharedReg727_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg727_out;
SharedReg728_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg728_out;
SharedReg729_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg729_out;
SharedReg730_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg730_out;
SharedReg831_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg831_out;
SharedReg92_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg92_out;
SharedReg656_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg656_out;
SharedReg742_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg742_out;
SharedReg833_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg833_out;
SharedReg779_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg779_out;
SharedReg497_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg497_out;
SharedReg789_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg789_out;
SharedReg651_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg651_out;
SharedReg835_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg835_out;
SharedReg822_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg822_out;
SharedReg823_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg823_out;
SharedReg824_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg824_out;
SharedReg825_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg825_out;
SharedReg826_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg826_out;
SharedReg827_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg827_out;
SharedReg752_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg760_out;
SharedReg789_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg789_out;
SharedReg715_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg715_out;
SharedReg762_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg762_out;
SharedReg470_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg470_out;
SharedReg805_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg805_out;
SharedReg719_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg719_out;
SharedReg861_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg861_out;
SharedReg216_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg216_out;
SharedReg92_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg92_out;
SharedReg722_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg722_out;
SharedReg815_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg815_out;
SharedReg672_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg672_out;
SharedReg218_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg218_out;
SharedReg770_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg770_out;
SharedReg771_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg771_out;
SharedReg718_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg718_out;
SharedReg809_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg809_out;
SharedReg720_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg720_out;
SharedReg842_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg842_out;
SharedReg816_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg816_out;
SharedReg496_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg496_out;
SharedReg814_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg814_out;
SharedReg693_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg693_out;
SharedReg724_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg725_out;
SharedReg847_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg847_out;
SharedReg235_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg235_out;
   MUX_Product11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg754_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg755_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg730_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg831_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg92_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg656_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg742_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg833_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg779_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg497_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg789_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg651_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg756_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg835_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg822_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg823_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg824_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg825_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg826_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg827_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg752_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg760_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg789_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg757_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg715_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg762_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg470_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg805_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg719_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg861_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg216_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg92_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg722_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg815_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg758_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg672_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg218_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg770_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg771_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg718_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg809_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg720_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg842_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg816_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg496_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg759_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg814_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg693_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg724_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg725_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg847_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg235_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg815_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg727_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg728_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg729_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product11_3_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_3_impl_0_out,
                 Y => Delay1No62_out);

SharedReg504_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg119_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg119_out;
SharedReg117_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg117_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg117_out;
SharedReg678_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg678_out;
SharedReg677_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg677_out;
SharedReg521_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg521_out;
SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg114_out;
SharedReg232_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg232_out;
SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg114_out;
SharedReg233_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg233_out;
SharedReg660_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg660_out;
SharedReg785_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg785_out;
SharedReg832_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg832_out;
SharedReg90_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg90_out;
SharedReg474_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg474_out;
SharedReg118_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg118_out;
SharedReg780_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg780_out;
SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg88_out;
SharedReg834_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg834_out;
SharedReg653_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg653_out;
SharedReg654_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg654_out;
SharedReg471_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg471_out;
SharedReg469_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg469_out;
SharedReg653_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg653_out;
SharedReg651_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg651_out;
SharedReg469_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg469_out;
SharedReg652_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg652_out;
SharedReg468_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg468_out;
SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg114_out;
SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg88_out;
SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg88_out;
SharedReg852_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg852_out;
SharedReg470_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg470_out;
SharedReg657_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg657_out;
SharedReg652_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg652_out;
SharedReg766_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg766_out;
SharedReg767_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg767_out;
SharedReg478_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg478_out;
SharedReg475_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg475_out;
SharedReg863_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg863_out;
SharedReg769_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg769_out;
SharedReg220_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg220_out;
SharedReg96_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg96_out;
SharedReg237_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg237_out;
SharedReg494_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg494_out;
SharedReg120_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg120_out;
SharedReg676_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg676_out;
SharedReg494_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg494_out;
SharedReg829_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg829_out;
SharedReg495_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg495_out;
SharedReg760_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg760_out;
SharedReg238_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg238_out;
SharedReg122_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg122_out;
SharedReg680_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg680_out;
SharedReg797_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg797_out;
   MUX_Product11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg119_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg233_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg660_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg785_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg832_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg90_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg474_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg118_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg780_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg834_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg117_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg653_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg654_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg471_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg469_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg653_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg651_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg469_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg652_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg468_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg117_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg88_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg852_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg470_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg657_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg652_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg766_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg767_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg478_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg475_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg678_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg863_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg769_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg220_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg96_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg237_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg494_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg120_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg676_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg494_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg829_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg677_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg495_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg760_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg238_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg122_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg680_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg797_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg521_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg232_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg114_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product11_3_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_3_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product11_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_4_impl_out,
                 X => Delay1No64_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg257_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg257_out;
SharedReg118_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
SharedReg114_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg114_out;
SharedReg494_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg494_out;
SharedReg673_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg673_out;
SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg672_out;
SharedReg677_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg677_out;
SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg672_out;
SharedReg698_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg698_out;
SharedReg674_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg674_out;
SharedReg816_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg816_out;
SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg672_out;
SharedReg718_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg718_out;
SharedReg720_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg720_out;
SharedReg804_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg804_out;
SharedReg809_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg809_out;
SharedReg842_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg842_out;
SharedReg843_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg843_out;
SharedReg858_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg858_out;
SharedReg727_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg727_out;
SharedReg729_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg729_out;
SharedReg742_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg742_out;
SharedReg717_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg717_out;
SharedReg728_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg728_out;
SharedReg778_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg778_out;
SharedReg850_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg850_out;
SharedReg724_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg724_out;
SharedReg853_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg853_out;
SharedReg768_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg768_out;
SharedReg831_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg831_out;
SharedReg833_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg833_out;
SharedReg757_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg757_out;
SharedReg756_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg756_out;
SharedReg751_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg751_out;
SharedReg750_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg750_out;
SharedReg841_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg841_out;
SharedReg748_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg748_out;
SharedReg749_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg749_out;
SharedReg838_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg838_out;
SharedReg725_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg725_out;
SharedReg758_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg758_out;
SharedReg747_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg747_out;
SharedReg822_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg822_out;
SharedReg754_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg754_out;
SharedReg752_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg752_out;
SharedReg755_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg755_out;
SharedReg753_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg753_out;
SharedReg822_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg822_out;
SharedReg835_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg835_out;
SharedReg716_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg716_out;
SharedReg862_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg862_out;
   MUX_Product11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_51_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg257_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg816_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg718_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg720_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg804_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg809_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg842_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg843_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg858_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg727_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg114_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg729_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg742_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg717_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg728_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg778_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg850_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg724_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg853_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg768_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg831_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg494_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg833_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg757_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg756_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg751_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg750_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg841_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg748_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg749_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg838_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg725_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg673_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg758_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg747_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg822_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg754_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg752_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg755_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg753_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg822_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg835_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg716_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg862_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_6 => SharedReg677_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg672_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg698_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg674_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product11_4_impl_0_LUT_out,
                 oMux => MUX_Product11_4_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_0_out,
                 Y => Delay1No64_out);

SharedReg259_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg146_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
SharedReg116_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg140_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg140_out;
SharedReg140_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg140_out;
SharedReg147_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
SharedReg254_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg254_out;
SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg143_out;
SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg143_out;
SharedReg141_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg141_out;
SharedReg254_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg254_out;
SharedReg141_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg141_out;
SharedReg256_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg256_out;
SharedReg115_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg115_out;
SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg143_out;
SharedReg145_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg145_out;
SharedReg257_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg257_out;
SharedReg146_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg146_out;
SharedReg260_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg260_out;
SharedReg148_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg148_out;
SharedReg232_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg232_out;
SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg517_out;
SharedReg694_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg694_out;
SharedReg514_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg514_out;
SharedReg497_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg497_out;
SharedReg681_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg681_out;
SharedReg527_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg527_out;
SharedReg701_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg701_out;
SharedReg518_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg518_out;
SharedReg492_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg492_out;
SharedReg492_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg492_out;
SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg517_out;
SharedReg693_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg693_out;
SharedReg675_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg675_out;
SharedReg674_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg674_out;
SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg517_out;
SharedReg697_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg697_out;
SharedReg700_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg700_out;
SharedReg701_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg701_out;
SharedReg693_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg693_out;
SharedReg763_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg763_out;
SharedReg761_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg761_out;
SharedReg785_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg785_out;
SharedReg832_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg832_out;
SharedReg840_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg840_out;
SharedReg839_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg839_out;
SharedReg803_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg803_out;
SharedReg837_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg837_out;
SharedReg796_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg796_out;
SharedReg834_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg834_out;
SharedReg760_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg760_out;
   MUX_Product11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_51_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg254_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg141_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg256_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg115_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg145_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg257_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg146_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg260_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg148_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg116_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg232_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg694_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg514_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg497_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg681_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg527_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg701_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg518_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg492_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg140_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg492_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg693_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg675_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg674_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg517_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg697_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg700_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg701_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg693_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg140_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg763_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg761_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg785_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg832_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg840_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg839_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg803_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg837_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg796_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg834_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg147_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg760_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_6 => SharedReg254_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg143_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg141_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product11_4_impl_1_LUT_out,
                 oMux => MUX_Product11_4_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No66_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg39_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg792_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg168_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg166_out;
SharedReg795_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg795_out;
SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg167_out;
SharedReg760_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg760_out;
SharedReg862_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg862_out;
SharedReg609_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg609_out;
SharedReg846_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg846_out;
SharedReg169_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg169_out;
SharedReg171_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg171_out;
SharedReg612_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg612_out;
SharedReg844_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg844_out;
SharedReg721_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg721_out;
SharedReg816_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg816_out;
SharedReg722_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg722_out;
SharedReg814_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg814_out;
SharedReg616_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg616_out;
SharedReg172_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg172_out;
SharedReg770_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg770_out;
SharedReg853_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg853_out;
SharedReg169_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg169_out;
SharedReg798_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg798_out;
SharedReg799_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg799_out;
SharedReg39_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg39_out;
SharedReg801_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg802_out;
SharedReg40_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg40_out;
SharedReg637_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg637_out;
SharedReg36_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg36_out;
SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg166_out;
SharedReg774_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg774_out;
SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg167_out;
SharedReg776_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg776_out;
SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg167_out;
SharedReg808_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg808_out;
SharedReg733_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg733_out;
SharedReg778_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg778_out;
SharedReg779_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg780_out;
SharedReg174_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg174_out;
SharedReg851_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg851_out;
SharedReg782_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg783_out;
SharedReg818_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg818_out;
SharedReg741_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg741_out;
SharedReg819_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg819_out;
SharedReg742_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg742_out;
SharedReg820_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg820_out;
SharedReg735_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg735_out;
SharedReg780_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg780_out;
SharedReg789_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg789_out;
SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg166_out;
SharedReg821_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg821_out;
SharedReg836_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg836_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg169_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg171_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg612_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg844_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg721_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg816_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg722_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg814_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg616_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg172_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg168_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg770_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg853_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg169_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg798_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg799_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg39_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg801_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg802_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg40_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg637_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg36_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg774_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg776_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg808_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg733_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg778_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg779_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg795_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg780_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg174_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg851_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg782_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg783_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg818_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg741_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg819_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg742_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg820_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg167_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg735_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg780_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg789_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg166_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg821_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg836_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg760_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg862_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg609_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg846_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No66_out);

SharedReg791_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg791_out;
SharedReg37_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg793_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg37_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg37_out;
SharedReg796_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg796_out;
SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg36_out;
SharedReg609_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg609_out;
SharedReg860_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg860_out;
SharedReg423_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg423_out;
SharedReg763_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg763_out;
SharedReg764_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg764_out;
SharedReg809_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg809_out;
SharedReg612_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg612_out;
SharedReg39_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg39_out;
SharedReg426_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg426_out;
SharedReg42_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg42_out;
SharedReg429_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg429_out;
SharedReg845_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg845_out;
SharedReg769_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg769_out;
SharedReg44_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg44_out;
SharedReg617_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg617_out;
SharedReg797_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg797_out;
SharedReg435_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg435_out;
SharedReg41_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg41_out;
SharedReg800_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg800_out;
SharedReg39_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg39_out;
SharedReg615_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg615_out;
SharedReg803_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg803_out;
SharedReg845_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg845_out;
SharedReg772_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg772_out;
SharedReg773_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg773_out;
SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg36_out;
SharedReg775_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg775_out;
SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg36_out;
SharedReg777_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg777_out;
SharedReg610_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg610_out;
SharedReg170_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg170_out;
SharedReg43_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg43_out;
SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg40_out;
SharedReg427_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg427_out;
SharedReg781_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg781_out;
SharedReg431_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg431_out;
SharedReg46_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg46_out;
SharedReg174_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg174_out;
SharedReg618_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg618_out;
SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg40_out;
SharedReg614_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg614_out;
SharedReg620_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg620_out;
SharedReg428_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg428_out;
SharedReg66_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg66_out;
SharedReg450_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg450_out;
SharedReg166_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg166_out;
SharedReg790_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg790_out;
SharedReg610_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg610_out;
SharedReg425_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg425_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg791_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg763_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg764_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg809_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg612_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg39_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg426_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg42_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg429_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg845_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg769_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg793_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg44_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg617_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg797_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg435_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg41_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg800_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg39_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg615_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg803_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg845_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg794_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg772_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg773_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg775_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg777_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg610_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg170_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg43_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg37_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg427_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg781_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg431_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg46_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg174_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg618_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg40_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg614_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg620_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg428_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg796_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg66_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg450_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg166_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg790_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg610_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg425_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg36_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg609_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg860_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg423_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product21_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_1_impl_out,
                 X => Delay1No68_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg818_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg818_out;
SharedReg741_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg741_out;
SharedReg819_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg819_out;
SharedReg742_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg742_out;
SharedReg820_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg820_out;
SharedReg735_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg735_out;
SharedReg780_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg780_out;
SharedReg789_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg789_out;
SharedReg188_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg188_out;
SharedReg821_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg821_out;
SharedReg836_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg836_out;
SharedReg65_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg65_out;
SharedReg792_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg792_out;
SharedReg190_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg190_out;
SharedReg188_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg188_out;
SharedReg795_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg795_out;
SharedReg189_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg189_out;
SharedReg760_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg760_out;
SharedReg862_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg862_out;
SharedReg630_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg630_out;
SharedReg846_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg846_out;
SharedReg191_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg191_out;
SharedReg193_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg193_out;
SharedReg633_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg633_out;
SharedReg844_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg844_out;
SharedReg721_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg721_out;
SharedReg816_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg816_out;
SharedReg722_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg722_out;
SharedReg814_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg814_out;
SharedReg862_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg862_out;
SharedReg194_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg194_out;
SharedReg770_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg770_out;
SharedReg853_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg853_out;
SharedReg753_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg753_out;
SharedReg754_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg758_out;
SharedReg759_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg759_out;
SharedReg723_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg723_out;
SharedReg727_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg727_out;
SharedReg848_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg848_out;
SharedReg806_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg806_out;
SharedReg630_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg630_out;
SharedReg811_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg811_out;
SharedReg807_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg807_out;
SharedReg631_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg631_out;
SharedReg849_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg849_out;
SharedReg637_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg637_out;
SharedReg92_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg92_out;
SharedReg723_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg723_out;
SharedReg737_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg737_out;
SharedReg857_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg857_out;
SharedReg817_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg817_out;
SharedReg453_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg453_out;
   MUX_Product21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg818_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg741_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg836_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg65_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg792_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg190_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg188_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg795_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg189_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg760_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg862_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg630_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg819_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg846_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg191_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg193_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg633_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg844_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg721_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg816_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg722_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg814_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg862_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg742_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg194_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg770_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg853_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg753_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg754_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg755_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg756_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg757_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg758_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg759_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg820_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg723_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg727_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg848_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg806_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg630_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg811_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg807_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg631_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg849_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg637_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg735_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg92_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg723_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg737_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg857_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg817_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg453_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg780_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg789_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg188_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg821_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product21_1_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_0_out,
                 Y => Delay1No68_out);

SharedReg639_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg639_out;
SharedReg66_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg635_out;
SharedReg641_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg641_out;
SharedReg451_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg451_out;
SharedReg92_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg92_out;
SharedReg473_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg473_out;
SharedReg188_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg188_out;
SharedReg790_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg790_out;
SharedReg631_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg631_out;
SharedReg448_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg448_out;
SharedReg791_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg791_out;
SharedReg63_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg63_out;
SharedReg793_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg794_out;
SharedReg63_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg63_out;
SharedReg796_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg796_out;
SharedReg62_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg62_out;
SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg630_out;
SharedReg860_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg860_out;
SharedReg446_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg446_out;
SharedReg763_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg763_out;
SharedReg764_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg764_out;
SharedReg809_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg809_out;
SharedReg633_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg633_out;
SharedReg65_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg65_out;
SharedReg449_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg449_out;
SharedReg68_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg68_out;
SharedReg452_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg452_out;
SharedReg651_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg651_out;
SharedReg769_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg769_out;
SharedReg70_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg70_out;
SharedReg638_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg638_out;
SharedReg77_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg77_out;
SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg635_out;
SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg635_out;
SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg635_out;
SharedReg191_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg191_out;
SharedReg449_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg449_out;
SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg635_out;
SharedReg216_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg216_out;
SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg630_out;
SharedReg445_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg445_out;
SharedReg445_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg445_out;
SharedReg855_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg855_out;
SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg630_out;
SharedReg631_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg631_out;
SharedReg812_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg812_out;
SharedReg634_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg634_out;
SharedReg856_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg856_out;
SharedReg803_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg803_out;
SharedReg238_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg238_out;
SharedReg451_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg451_out;
SharedReg454_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg454_out;
SharedReg452_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg452_out;
SharedReg830_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg830_out;
   MUX_Product21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg639_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg448_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg791_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg63_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg793_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg794_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg63_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg796_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg62_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg860_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg446_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg763_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg764_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg809_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg633_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg65_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg449_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg68_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg452_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg651_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg641_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg769_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg70_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg638_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg77_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg191_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg449_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg635_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg451_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg216_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg445_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg445_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg855_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg630_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg631_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg812_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg634_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg856_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg92_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg803_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg238_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg451_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg454_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg452_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg830_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg473_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg188_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg790_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg631_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product21_1_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product21_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_2_impl_out,
                 X => Delay1No70_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg811_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg811_out;
SharedReg807_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg652_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg652_out;
SharedReg849_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg849_out;
SharedReg658_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg658_out;
SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg118_out;
SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg814_out;
SharedReg737_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg737_out;
SharedReg857_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg857_out;
SharedReg817_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg817_out;
SharedReg476_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg476_out;
SharedReg818_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg818_out;
SharedReg741_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg741_out;
SharedReg819_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg819_out;
SharedReg742_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg742_out;
SharedReg820_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg820_out;
SharedReg735_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg735_out;
SharedReg780_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg780_out;
SharedReg789_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg789_out;
SharedReg210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg210_out;
SharedReg821_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg821_out;
SharedReg836_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg836_out;
SharedReg91_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg91_out;
SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg792_out;
SharedReg212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg212_out;
SharedReg210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg210_out;
SharedReg795_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg795_out;
SharedReg211_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg211_out;
SharedReg760_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg760_out;
SharedReg789_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg789_out;
SharedReg651_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg651_out;
SharedReg846_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg846_out;
SharedReg213_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg213_out;
SharedReg718_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg718_out;
SharedReg213_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg213_out;
SharedReg859_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg859_out;
SharedReg766_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg766_out;
SharedReg828_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg828_out;
SharedReg768_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg768_out;
SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg814_out;
SharedReg863_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg863_out;
SharedReg724_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg725_out;
SharedReg726_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg726_out;
SharedReg797_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg797_out;
SharedReg656_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg656_out;
SharedReg799_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg799_out;
SharedReg656_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg656_out;
SharedReg801_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg802_out;
SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg814_out;
SharedReg760_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg760_out;
SharedReg651_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg651_out;
SharedReg854_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg854_out;
SharedReg810_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg810_out;
SharedReg753_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg753_out;
   MUX_Product21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg811_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg476_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg818_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg741_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg819_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg742_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg820_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg735_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg780_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg789_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg652_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg821_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg836_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg91_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg212_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg210_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg795_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg211_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg760_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg789_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg651_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg846_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg213_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg718_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg213_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg859_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg766_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg828_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg768_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg658_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg863_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg724_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg725_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg726_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg797_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg656_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg799_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg656_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg801_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg802_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg118_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg760_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg651_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg854_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg810_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg753_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg814_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg737_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg857_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg817_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product21_2_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_0_out,
                 Y => Delay1No70_out);

SharedReg651_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg651_out;
SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg652_out;
SharedReg812_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg812_out;
SharedReg655_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg655_out;
SharedReg856_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg856_out;
SharedReg803_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg803_out;
SharedReg518_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg518_out;
SharedReg474_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg474_out;
SharedReg477_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg477_out;
SharedReg475_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg475_out;
SharedReg830_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg830_out;
SharedReg660_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg660_out;
SharedReg92_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg92_out;
SharedReg656_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg656_out;
SharedReg662_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg662_out;
SharedReg474_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg474_out;
SharedReg118_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg118_out;
SharedReg496_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg496_out;
SharedReg210_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg210_out;
SharedReg790_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg790_out;
SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg652_out;
SharedReg471_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg471_out;
SharedReg791_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg791_out;
SharedReg89_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg89_out;
SharedReg793_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg794_out;
SharedReg89_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg89_out;
SharedReg796_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg796_out;
SharedReg88_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg88_out;
SharedReg232_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg232_out;
SharedReg860_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg860_out;
SharedReg469_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg469_out;
SharedReg763_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg763_out;
SharedReg214_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg214_out;
SharedReg765_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg765_out;
SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg652_out;
SharedReg212_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg212_out;
SharedReg471_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg471_out;
SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg94_out;
SharedReg472_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg472_out;
SharedReg491_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg491_out;
SharedReg218_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg218_out;
SharedReg220_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg220_out;
SharedReg96_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg96_out;
SharedReg103_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg103_out;
SharedReg798_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg798_out;
SharedReg656_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg656_out;
SharedReg800_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg800_out;
SharedReg213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg213_out;
SharedReg472_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg472_out;
SharedReg498_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg498_out;
SharedReg514_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg514_out;
SharedReg772_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg772_out;
SharedReg468_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg468_out;
SharedReg468_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg468_out;
SharedReg235_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg235_out;
   MUX_Product21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg651_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg830_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg660_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg92_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg656_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg662_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg474_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg118_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg496_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg210_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg790_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg812_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg471_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg791_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg89_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg793_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg794_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg89_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg796_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg88_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg232_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg655_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg860_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg469_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg763_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg214_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg765_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg652_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg212_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg471_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg94_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg472_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg856_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg491_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg218_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg220_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg96_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg103_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg798_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg656_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg800_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg213_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg472_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg803_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg498_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg514_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg772_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg468_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg468_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg235_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg518_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg474_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg477_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg475_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product21_2_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product21_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_3_impl_out,
                 X => Delay1No72_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg235_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg235_out;
SharedReg126_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg126_out;
SharedReg240_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg240_out;
SharedReg233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg233_out;
SharedReg232_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg232_out;
SharedReg144_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg144_out;
SharedReg234_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg234_out;
SharedReg117_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg117_out;
SharedReg235_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg235_out;
SharedReg233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg233_out;
SharedReg672_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg672_out;
SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg828_out;
SharedReg519_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg519_out;
SharedReg672_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg672_out;
SharedReg760_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg760_out;
SharedReg718_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg718_out;
SharedReg851_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg851_out;
SharedReg859_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg859_out;
SharedReg735_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg735_out;
SharedReg776_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg776_out;
SharedReg741_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg741_out;
SharedReg784_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg784_out;
SharedReg743_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg743_out;
SharedReg783_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg783_out;
SharedReg778_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg778_out;
SharedReg727_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg727_out;
SharedReg786_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg786_out;
SharedReg806_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg806_out;
SharedReg787_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg787_out;
SharedReg733_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg733_out;
SharedReg782_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg782_out;
SharedReg780_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg780_out;
SharedReg808_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg808_out;
SharedReg848_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg848_out;
SharedReg846_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg846_out;
SharedReg768_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg768_out;
SharedReg795_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg795_out;
SharedReg757_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg757_out;
SharedReg792_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg792_out;
SharedReg758_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg758_out;
SharedReg752_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg752_out;
SharedReg797_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg797_out;
SharedReg758_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg758_out;
SharedReg756_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg756_out;
SharedReg822_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg822_out;
SharedReg746_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg746_out;
SharedReg745_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg745_out;
SharedReg755_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg755_out;
SharedReg754_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg754_out;
SharedReg725_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg725_out;
SharedReg724_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg724_out;
SharedReg726_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg726_out;
SharedReg766_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg766_out;
   MUX_Product21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_53_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg672_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg519_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg672_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg760_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg718_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg851_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg859_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg735_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg776_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg240_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg741_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg784_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg743_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg783_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg778_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg727_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg786_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg806_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg787_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg733_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg782_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg780_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg808_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg848_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg846_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg768_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg795_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg757_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg792_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg758_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg232_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg752_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg797_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg758_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg756_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg822_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg746_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg745_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg755_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg754_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg725_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg144_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg724_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg726_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg766_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_6 => SharedReg234_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg117_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg235_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg233_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product21_3_impl_0_LUT_out,
                 oMux => MUX_Product21_3_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_0_out,
                 Y => Delay1No72_out);

SharedReg236_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg236_out;
SharedReg114_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg114_out;
SharedReg116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg124_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg124_out;
SharedReg236_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg236_out;
SharedReg123_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg122_out;
SharedReg240_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg240_out;
SharedReg121_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg121_out;
SharedReg115_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg115_out;
SharedReg235_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg235_out;
SharedReg115_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg115_out;
SharedReg129_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg129_out;
SharedReg255_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg255_out;
SharedReg234_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg234_out;
SharedReg116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg116_out;
SharedReg232_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg232_out;
SharedReg120_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg120_out;
SharedReg242_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg242_out;
SharedReg240_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg240_out;
SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg122_out;
SharedReg144_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg144_out;
SharedReg114_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg114_out;
SharedReg494_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg494_out;
SharedReg500_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg500_out;
SharedReg682_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg682_out;
SharedReg672_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg672_out;
SharedReg491_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg491_out;
SharedReg491_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg491_out;
SharedReg495_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg495_out;
SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg677_out;
SharedReg699_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg699_out;
SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg677_out;
SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg677_out;
SharedReg673_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg673_out;
SharedReg494_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg494_out;
SharedReg492_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg492_out;
SharedReg829_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg829_out;
SharedReg519_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg519_out;
SharedReg673_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg673_out;
SharedReg763_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg763_out;
SharedReg855_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg855_out;
SharedReg860_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg860_out;
SharedReg777_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg777_out;
SharedReg788_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg788_out;
SharedReg781_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg781_out;
SharedReg794_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg794_out;
SharedReg803_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg803_out;
SharedReg793_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg793_out;
SharedReg796_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg796_out;
SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg791_out;
SharedReg765_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg765_out;
   MUX_Product21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_53_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg236_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg115_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg235_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg115_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg129_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg255_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg234_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg232_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg120_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg242_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg116_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg240_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg144_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg114_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg494_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg500_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg682_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg672_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg491_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg491_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg127_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg495_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg699_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg677_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg673_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg494_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg492_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg829_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg519_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg124_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg673_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg763_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg855_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg860_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg777_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg788_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg781_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg794_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg803_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg793_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg236_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg796_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg791_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg765_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_6 => SharedReg123_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg240_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg121_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product21_3_impl_1_LUT_out,
                 oMux => MUX_Product21_3_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product31_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_4_impl_out,
                 X => Delay1No74_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast);

SharedReg259_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg152_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg140_out;
SharedReg254_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg254_out;
SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg143_out;
SharedReg254_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg254_out;
SharedReg256_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg256_out;
SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg143_out;
SharedReg257_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg257_out;
SharedReg260_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg260_out;
SharedReg260_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg260_out;
SharedReg694_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg694_out;
SharedReg698_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg698_out;
SharedReg700_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg700_out;
SharedReg696_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg696_out;
SharedReg816_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg816_out;
SharedReg700_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg700_out;
SharedReg516_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg516_out;
SharedReg693_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg693_out;
SharedReg844_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg844_out;
SharedReg738_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg738_out;
SharedReg731_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg731_out;
SharedReg732_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg732_out;
SharedReg741_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg741_out;
SharedReg784_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg784_out;
SharedReg730_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg730_out;
SharedReg774_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg774_out;
SharedReg740_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg740_out;
SharedReg786_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg786_out;
SharedReg808_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg808_out;
SharedReg743_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg743_out;
SharedReg787_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg787_out;
SharedReg739_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg739_out;
SharedReg846_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg846_out;
SharedReg801_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg801_out;
SharedReg795_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg795_out;
SharedReg792_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg792_out;
SharedReg721_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg721_out;
SharedReg770_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg770_out;
SharedReg802_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg802_out;
SharedReg744_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg744_out;
SharedReg836_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg836_out;
SharedReg798_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg798_out;
SharedReg799_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg799_out;
SharedReg746_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg746_out;
SharedReg745_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg745_out;
SharedReg726_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg726_out;
SharedReg722_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg722_out;
SharedReg862_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg862_out;
   MUX_Product31_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_49_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg260_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg694_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg698_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg700_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg696_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg816_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg700_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg516_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg693_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg844_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg140_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg738_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg731_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg732_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg741_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg784_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg730_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg774_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg740_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg786_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg808_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg254_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg743_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg787_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg739_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg846_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg801_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg795_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg792_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg721_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg770_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg802_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg744_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg836_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg798_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg799_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg746_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg745_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg726_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg722_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg862_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_5 => SharedReg254_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg256_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg143_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg257_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg260_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product31_4_impl_0_LUT_out,
                 oMux => MUX_Product31_4_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_0_out,
                 Y => Delay1No74_out);

SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg153_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg153_out;
SharedReg150_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg150_out;
SharedReg149_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg149_out;
SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg148_out;
SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg140_out;
SharedReg255_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg255_out;
SharedReg262_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg262_out;
SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg143_out;
SharedReg141_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg141_out;
SharedReg141_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg141_out;
SharedReg254_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg254_out;
SharedReg145_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg145_out;
SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg142_out;
SharedReg254_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg254_out;
SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg148_out;
SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg143_out;
SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg148_out;
SharedReg261_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg261_out;
SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg140_out;
SharedReg255_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg255_out;
SharedReg517_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg517_out;
SharedReg527_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg527_out;
SharedReg524_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg524_out;
SharedReg693_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg693_out;
SharedReg703_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg703_out;
SharedReg697_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg697_out;
SharedReg518_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg518_out;
SharedReg518_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg518_out;
SharedReg696_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg696_out;
SharedReg515_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg515_out;
SharedReg764_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg764_out;
SharedReg809_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg809_out;
SharedReg845_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg845_out;
SharedReg860_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg860_out;
SharedReg781_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg781_out;
SharedReg772_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg772_out;
SharedReg773_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg773_out;
SharedReg813_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg813_out;
SharedReg788_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg788_out;
SharedReg856_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg856_out;
SharedReg852_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg852_out;
SharedReg769_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg769_out;
SharedReg800_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg800_out;
SharedReg794_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg794_out;
SharedReg793_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg793_out;
SharedReg791_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg791_out;
SharedReg796_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg796_out;
SharedReg797_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg797_out;
   MUX_Product31_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_49_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg141_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg254_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg145_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg142_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg254_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg261_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg150_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg255_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg517_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg527_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg524_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg693_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg703_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg697_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg518_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg518_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg696_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg149_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg515_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg764_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg809_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg845_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg860_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg781_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg772_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg773_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg813_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg788_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg148_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg856_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg852_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg769_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg800_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg794_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg793_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg791_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg796_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg797_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_5 => SharedReg140_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg255_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg262_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg143_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg141_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product31_4_impl_1_LUT_out,
                 oMux => MUX_Product31_4_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No76_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg180_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg180_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg283_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg283_out;
SharedReg285_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg285_out;
SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg282_out;
SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg280_out;
SharedReg542_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg542_out;
SharedReg586_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg586_out;
SharedReg281_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg281_out;
SharedReg587_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg587_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg276_out;
SharedReg438_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg438_out;
SharedReg441_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg441_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg277_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg358_out;
SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg280_out;
SharedReg361_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg361_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg276_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg276_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg422_out;
SharedReg620_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg620_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg422_out;
SharedReg45_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg45_out;
SharedReg432_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg432_out;
SharedReg48_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg48_out;
SharedReg544_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg544_out;
SharedReg544_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg544_out;
SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg282_out;
SharedReg281_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg281_out;
SharedReg543_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg543_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg277_out;
SharedReg435_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg435_out;
SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg277_out;
SharedReg538_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg538_out;
SharedReg542_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg542_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg276_out;
SharedReg426_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg426_out;
SharedReg614_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg614_out;
SharedReg278_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg278_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg358_out;
SharedReg427_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg427_out;
SharedReg172_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg172_out;
SharedReg278_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg278_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg276_out;
SharedReg428_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg428_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg358_out;
SharedReg538_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg538_out;
SharedReg432_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg432_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg422_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg180_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg285_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg542_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg586_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg281_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg587_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg438_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg441_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg2_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg280_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg361_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg620_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg45_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg14_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg432_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg48_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg544_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg544_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg281_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg543_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg435_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg277_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg4_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg538_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg542_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg426_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg614_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg278_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg427_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg172_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg278_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg7_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg276_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg428_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg358_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg538_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg432_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg422_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg10_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg283_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No76_out);

SharedReg186_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg366_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg366_out;
SharedReg364_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg364_out;
SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg363_out;
SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg363_out;
SharedReg591_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg591_out;
SharedReg588_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg588_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg358_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg358_out;
SharedReg361_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg361_out;
SharedReg434_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg434_out;
SharedReg444_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg444_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg276_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg276_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg358_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg358_out;
SharedReg590_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg590_out;
SharedReg547_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg547_out;
SharedReg613_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg613_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg422_out;
SharedReg610_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg610_out;
SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg36_out;
SharedReg423_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg423_out;
SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg167_out;
SharedReg548_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg548_out;
Delay25No20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast <= Delay25No20_out;
SharedReg366_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg366_out;
SharedReg364_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg364_out;
SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg362_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg358_out;
SharedReg423_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg423_out;
SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg358_out;
SharedReg537_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg537_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg276_out;
SharedReg365_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg365_out;
SharedReg440_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg440_out;
SharedReg627_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg627_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg276_out;
SharedReg546_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg546_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg422_out;
SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg167_out;
SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg362_out;
SharedReg368_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg368_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg422_out;
SharedReg597_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg597_out;
SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg276_out;
SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg422_out;
SharedReg609_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg609_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg364_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg591_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg588_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg361_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg434_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg444_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg590_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg547_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg613_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg610_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg36_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg32_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg423_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg548_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay25No20_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg366_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg364_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg423_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg358_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg537_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg365_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg440_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg627_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg546_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg362_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg368_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg597_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg276_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg422_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg609_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg28_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg27_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg366_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No78_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg360_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg360_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg287_out;
SharedReg450_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg450_out;
SharedReg194_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg194_out;
SharedReg588_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg588_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg287_out;
SharedReg451_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg451_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg370_out;
SharedReg551_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg551_out;
SharedReg455_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg455_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg445_out;
SharedReg202_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg202_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg8_out;
SharedReg294_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg294_out;
SharedReg296_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg296_out;
SharedReg293_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg293_out;
SharedReg291_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg291_out;
SharedReg554_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg554_out;
SharedReg322_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg322_out;
SharedReg292_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg292_out;
SharedReg323_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg323_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg287_out;
SharedReg461_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg461_out;
SharedReg464_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg464_out;
SharedReg288_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg288_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg370_out;
SharedReg291_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg291_out;
SharedReg373_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg373_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg287_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg287_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg445_out;
SharedReg641_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg641_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg445_out;
SharedReg71_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg71_out;
SharedReg455_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg455_out;
SharedReg74_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg74_out;
SharedReg556_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg556_out;
SharedReg377_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg377_out;
SharedReg591_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg591_out;
SharedReg590_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg590_out;
SharedReg376_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg376_out;
SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg587_out;
SharedReg458_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg458_out;
SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg587_out;
SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg371_out;
SharedReg375_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg375_out;
SharedReg586_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg586_out;
SharedReg449_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg449_out;
SharedReg635_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg635_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg360_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg202_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg2_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg14_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg4_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg7_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg10_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg9_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg8_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg450_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg294_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg296_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg293_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg291_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg554_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg322_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg292_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg323_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg461_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg194_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg464_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg288_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg291_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg373_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg641_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg445_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg588_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg71_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg455_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg74_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg556_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg377_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg591_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg590_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg376_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg458_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg587_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg371_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg375_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg586_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg449_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg635_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg451_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg370_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg551_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg455_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No78_out);

SharedReg586_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg586_out;
SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg379_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg445_out;
SharedReg189_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg189_out;
SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg291_out;
SharedReg297_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg297_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg445_out;
SharedReg562_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg287_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg630_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg630_out;
SharedReg208_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg208_out;
SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg26_out;
SharedReg378_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg378_out;
SharedReg376_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg376_out;
SharedReg375_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg375_out;
SharedReg375_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg375_out;
SharedReg327_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg327_out;
SharedReg324_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg324_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg370_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg370_out;
SharedReg373_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg373_out;
SharedReg457_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg457_out;
SharedReg467_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg467_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg287_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg287_out;
SharedReg358_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg358_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg370_out;
SharedReg326_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg326_out;
SharedReg559_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg559_out;
SharedReg634_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg634_out;
SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg445_out;
SharedReg631_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg631_out;
SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg62_out;
SharedReg446_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg446_out;
SharedReg189_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg189_out;
SharedReg561_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg561_out;
Delay25No21_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast <= Delay25No21_out;
SharedReg295_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg295_out;
SharedReg293_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg293_out;
SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg291_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg287_out;
SharedReg446_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg446_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg287_out;
SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg370_out;
SharedReg586_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg586_out;
SharedReg294_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg294_out;
SharedReg463_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg463_out;
SharedReg648_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg648_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg586_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg630_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg208_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg18_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg20_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg32_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg25_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg28_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg27_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg378_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg376_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg375_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg375_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg327_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg324_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg373_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg457_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg189_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg467_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg358_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg326_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg559_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg634_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg631_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg62_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg446_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg189_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg561_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => Delay25No21_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg295_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg293_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg291_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg446_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg297_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg370_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg586_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg294_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg463_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg648_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg287_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No80_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg555_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg555_out;
SharedReg554_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg554_out;
SharedReg304_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg304_out;
SharedReg551_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg551_out;
SharedReg481_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg481_out;
SharedReg323_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg323_out;
SharedReg384_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg384_out;
SharedReg303_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg303_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg322_out;
SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg472_out;
SharedReg656_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg656_out;
SharedReg372_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg372_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg298_out;
SharedReg473_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg473_out;
SharedReg216_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg216_out;
SharedReg324_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg324_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg298_out;
SharedReg474_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg474_out;
SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg383_out;
SharedReg334_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg334_out;
SharedReg478_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg478_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg468_out;
SharedReg224_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg224_out;
SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg8_out;
SharedReg305_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg305_out;
SharedReg308_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg308_out;
SharedReg304_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg304_out;
SharedReg302_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg302_out;
SharedReg337_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg337_out;
SharedReg310_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg310_out;
SharedReg303_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg303_out;
SharedReg334_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg334_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg322_out;
SharedReg484_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg484_out;
SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg487_out;
SharedReg323_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg323_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg298_out;
SharedReg325_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg325_out;
SharedReg301_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg301_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg322_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg322_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg468_out;
SharedReg662_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg662_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg468_out;
SharedReg97_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg97_out;
SharedReg478_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg478_out;
SharedReg100_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg100_out;
SharedReg390_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg390_out;
SharedReg305_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg305_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg555_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg554_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg656_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg372_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg473_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg216_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg324_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg474_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg334_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg304_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg478_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg224_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg2_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg14_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg4_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg7_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg10_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg9_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg551_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg8_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg305_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg308_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg304_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg302_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg337_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg310_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg303_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg334_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg481_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg484_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg487_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg323_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg298_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg325_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg301_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg662_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg323_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg468_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg97_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg478_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg100_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg390_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg305_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg384_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg303_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg322_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg472_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No80_out);

SharedReg329_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg329_out;
SharedReg327_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg327_out;
SharedReg374_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg374_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg322_out;
SharedReg469_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg469_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg298_out;
SharedReg383_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg383_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg322_out;
SharedReg328_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg328_out;
SharedReg486_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg486_out;
SharedReg669_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg669_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg322_out;
SharedReg307_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg307_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg468_out;
SharedReg211_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg211_out;
SharedReg302_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg302_out;
SharedReg332_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg332_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg468_out;
SharedReg394_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg394_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg298_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg468_out;
SharedReg651_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg651_out;
SharedReg230_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg230_out;
SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg26_out;
SharedReg391_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg389_out;
SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg388_out;
SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg388_out;
SharedReg316_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg316_out;
SharedReg312_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg312_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg298_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg298_out;
SharedReg386_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg386_out;
SharedReg480_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg480_out;
SharedReg490_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg490_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg322_out;
SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg322_out;
SharedReg287_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg287_out;
SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg298_out;
SharedReg337_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg337_out;
SharedReg343_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg343_out;
SharedReg655_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg655_out;
SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg468_out;
SharedReg652_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg652_out;
SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg88_out;
SharedReg469_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg469_out;
SharedReg211_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg211_out;
SharedReg393_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg393_out;
Delay25No22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast <= Delay25No22_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg329_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg669_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg307_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg211_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg302_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg332_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg394_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg374_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg651_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg230_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg18_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg20_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg32_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg25_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg28_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg26_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg391_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg389_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg388_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg316_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg312_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg386_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg469_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg480_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg490_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg287_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg337_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg343_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg655_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg468_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg298_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg652_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg88_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg469_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg211_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg393_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => Delay25No22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg383_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg322_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg328_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg486_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No82_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg313_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg313_out;
SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg333_out;
SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg333_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg491_out;
SharedReg683_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg683_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg491_out;
SharedReg123_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg123_out;
SharedReg501_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg501_out;
SharedReg126_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg126_out;
SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg403_out;
SharedReg317_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg317_out;
SharedReg338_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg338_out;
SharedReg337_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg337_out;
SharedReg402_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg402_out;
SharedReg334_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg334_out;
SharedReg504_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg504_out;
SharedReg311_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg311_out;
SharedReg575_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg575_out;
SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg401_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg310_out;
SharedReg495_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg495_out;
SharedReg677_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg677_out;
SharedReg385_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg385_out;
SharedReg396_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg396_out;
SharedReg496_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg496_out;
SharedReg238_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg238_out;
SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg312_out;
SharedReg396_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg396_out;
SharedReg497_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg497_out;
SharedReg574_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg574_out;
SharedReg346_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg346_out;
SharedReg501_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg501_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg491_out;
SharedReg246_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg246_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg8_out;
SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg403_out;
SharedReg308_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg308_out;
SharedReg316_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg316_out;
SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg314_out;
SharedReg579_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg579_out;
SharedReg345_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg345_out;
SharedReg315_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg315_out;
SharedReg575_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg575_out;
SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg333_out;
SharedReg507_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg507_out;
SharedReg510_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg510_out;
SharedReg334_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg334_out;
SharedReg383_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg383_out;
SharedReg336_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg336_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg313_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg317_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg338_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg337_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg402_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg334_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg504_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg311_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg575_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg401_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg310_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg495_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg677_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg385_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg396_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg496_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg238_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg396_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg497_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg574_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg346_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg501_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg246_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg2_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg14_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg4_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg7_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg10_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg683_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg9_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg8_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg308_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg316_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg579_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg345_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg315_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg575_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg491_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg333_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg507_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg510_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg334_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg383_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg336_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg123_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg501_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg126_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No82_out);

SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg310_out;
SharedReg579_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg579_out;
SharedReg583_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg583_out;
SharedReg676_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg676_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg491_out;
SharedReg673_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg673_out;
SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg114_out;
SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg492_out;
SharedReg233_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg233_out;
SharedReg406_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg406_out;
SharedReg409_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg409_out;
SharedReg340_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg340_out;
SharedReg316_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg316_out;
SharedReg387_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg387_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg310_out;
SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg492_out;
SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg396_out;
SharedReg574_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg574_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg310_out;
SharedReg317_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg317_out;
SharedReg509_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg509_out;
SharedReg690_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg690_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg310_out;
SharedReg405_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg405_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg491_out;
SharedReg233_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg233_out;
SharedReg400_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg400_out;
SharedReg320_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg320_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg491_out;
SharedReg584_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg584_out;
SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg396_out;
SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg491_out;
SharedReg672_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg672_out;
SharedReg252_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg252_out;
SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg26_out;
SharedReg582_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg582_out;
SharedReg402_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg402_out;
SharedReg401_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg401_out;
SharedReg401_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg401_out;
SharedReg351_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg351_out;
SharedReg347_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg347_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg310_out;
SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg310_out;
SharedReg399_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg399_out;
SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg503_out;
SharedReg513_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg513_out;
SharedReg333_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg333_out;
SharedReg298_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg298_out;
SharedReg287_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg287_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg579_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg409_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg340_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg316_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg387_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg574_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg317_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg583_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg509_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg690_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg405_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg233_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg400_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg320_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg584_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg676_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg396_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg672_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg252_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg18_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg20_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg32_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg25_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg491_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg27_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg26_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg582_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg402_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg401_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg401_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg351_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg347_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg310_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg673_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg399_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg503_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg513_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg333_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg298_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg287_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg114_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg492_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg233_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg406_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No84_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg351_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg349_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg349_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg568_out;
SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg563_out;
SharedReg326_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg599_out;
SharedReg345_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg345_out;
SharedReg530_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg530_out;
SharedReg533_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg533_out;
SharedReg346_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg346_out;
SharedReg298_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg298_out;
SharedReg349_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg349_out;
SharedReg577_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg577_out;
SharedReg345_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg345_out;
SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg574_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg514_out;
SharedReg704_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg704_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg514_out;
SharedReg149_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg149_out;
SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg524_out;
SharedReg152_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg152_out;
SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg416_out;
SharedReg570_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg570_out;
SharedReg351_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg351_out;
SharedReg350_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg350_out;
SharedReg569_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg569_out;
SharedReg346_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg346_out;
SharedReg527_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg527_out;
SharedReg411_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg411_out;
SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg599_out;
SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg568_out;
SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg574_out;
SharedReg518_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg518_out;
SharedReg698_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg698_out;
SharedReg398_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg398_out;
SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg563_out;
SharedReg519_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg519_out;
SharedReg260_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg260_out;
SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg412_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg410_out;
SharedReg520_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg520_out;
SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg563_out;
SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg599_out;
SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg524_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg514_out;
SharedReg268_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg268_out;
SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg_out;
SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg2_out;
SharedReg14_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg14_out;
SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg4_out;
SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg7_out;
SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg10_out;
SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg9_out;
SharedReg8_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg8_out;
SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg416_out;
SharedReg418_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg418_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg349_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg298_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg349_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg577_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg345_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg704_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg149_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg152_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg570_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg351_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg350_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg569_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg346_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg527_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg411_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg568_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg574_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg518_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg698_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg398_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg519_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg260_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg412_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg410_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg326_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg520_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg563_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg524_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg514_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg268_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg2_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg14_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg4_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg599_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg7_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg10_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg9_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg8_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg416_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg418_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg345_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg530_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg533_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg346_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No84_out);

SharedReg414_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg414_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg414_out;
SharedReg604_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg604_out;
SharedReg600_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg600_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg410_out;
SharedReg348_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg348_out;
SharedReg526_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg526_out;
SharedReg536_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg536_out;
SharedReg396_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg396_out;
SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg322_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg410_out;
SharedReg603_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg603_out;
SharedReg419_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg419_out;
SharedReg697_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg697_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg514_out;
SharedReg694_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg694_out;
SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg140_out;
SharedReg515_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg515_out;
SharedReg255_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg255_out;
SharedReg573_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg573_out;
SharedReg585_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg585_out;
SharedReg417_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg417_out;
SharedReg415_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg415_out;
SharedReg400_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg400_out;
SharedReg563_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg563_out;
SharedReg515_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg515_out;
SharedReg563_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg563_out;
SharedReg598_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg598_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg410_out;
SharedReg416_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg416_out;
SharedReg532_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg532_out;
SharedReg711_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg711_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg410_out;
SharedReg607_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg607_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg514_out;
SharedReg255_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg255_out;
SharedReg567_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg567_out;
SharedReg420_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg420_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg514_out;
Delay19No19_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast <= Delay19No19_out;
SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg410_out;
SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg514_out;
SharedReg693_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg693_out;
SharedReg274_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg274_out;
SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg20_out;
SharedReg32_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg32_out;
SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg22_out;
SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg25_out;
SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg28_out;
SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg27_out;
SharedReg26_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg26_out;
SharedReg571_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg571_out;
SharedReg415_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg415_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg414_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg603_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg419_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg697_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg694_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg140_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg515_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg604_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg255_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg573_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg585_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg417_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg415_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg400_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg563_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg515_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg563_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg598_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg600_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg416_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg532_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg711_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg607_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg255_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg567_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg420_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => Delay19No19_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg514_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg693_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg274_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg18_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg20_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg32_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg410_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg25_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg28_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg27_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg26_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg571_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg415_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg348_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg526_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg536_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg396_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Product12_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_0_impl_out,
                 X => Delay1No86_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg823_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg823_out;
SharedReg824_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg824_out;
SharedReg825_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg825_out;
SharedReg826_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg826_out;
SharedReg827_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg827_out;
SharedReg752_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg760_out;
SharedReg863_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg863_out;
SharedReg715_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg715_out;
SharedReg762_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg762_out;
SharedReg424_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg424_out;
SharedReg718_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg718_out;
SharedReg169_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg169_out;
SharedReg859_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg859_out;
SharedReg766_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg766_out;
SharedReg828_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg828_out;
SharedReg768_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg768_out;
SharedReg814_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg814_out;
SharedReg723_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg723_out;
SharedReg724_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg725_out;
SharedReg726_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg726_out;
SharedReg753_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg753_out;
SharedReg754_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg758_out;
SharedReg759_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg759_out;
SharedReg723_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg723_out;
SharedReg727_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg727_out;
SharedReg848_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg848_out;
SharedReg806_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg806_out;
SharedReg609_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg609_out;
SharedReg811_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg811_out;
SharedReg807_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg807_out;
SharedReg610_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg610_out;
SharedReg849_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg849_out;
SharedReg616_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg616_out;
SharedReg850_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg850_out;
SharedReg428_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg428_out;
SharedReg737_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg737_out;
SharedReg857_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg857_out;
SharedReg817_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg817_out;
SharedReg430_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg430_out;
SharedReg831_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg831_out;
SharedReg40_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg40_out;
SharedReg614_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg614_out;
SharedReg742_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg742_out;
SharedReg833_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg833_out;
SharedReg779_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg779_out;
SharedReg451_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg451_out;
SharedReg789_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg789_out;
SharedReg609_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg609_out;
SharedReg835_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg835_out;
SharedReg822_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg822_out;
   MUX_Product12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg823_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg824_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg424_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg718_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg169_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg859_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg766_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg828_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg768_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg814_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg723_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg724_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg825_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg725_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg726_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg753_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg754_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg755_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg756_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg757_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg758_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg759_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg723_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg826_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg727_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg848_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg806_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg609_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg811_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg807_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg610_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg849_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg616_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg850_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg827_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg428_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg737_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg857_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg817_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg430_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg831_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg40_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg614_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg742_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg833_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg752_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg779_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg451_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg789_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg609_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg835_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg822_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg760_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg863_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg715_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg762_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product12_0_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_0_out,
                 Y => Delay1No86_out);

SharedReg425_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg425_out;
SharedReg423_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg423_out;
SharedReg611_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg611_out;
SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg609_out;
SharedReg423_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg610_out;
SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg422_out;
SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg36_out;
SharedReg852_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg852_out;
SharedReg170_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg170_out;
SharedReg765_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg765_out;
SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg610_out;
SharedReg168_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg168_out;
SharedReg425_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg425_out;
SharedReg42_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg42_out;
SharedReg426_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg426_out;
SharedReg172_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg172_out;
SharedReg174_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg174_out;
SharedReg176_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg176_out;
SharedReg44_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg44_out;
SharedReg51_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg51_out;
SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg614_out;
SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg614_out;
SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg614_out;
SharedReg169_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg169_out;
SharedReg426_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg426_out;
SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg614_out;
SharedReg194_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg194_out;
SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg609_out;
SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg422_out;
SharedReg855_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg855_out;
SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg609_out;
SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg610_out;
SharedReg812_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg812_out;
SharedReg613_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg613_out;
SharedReg856_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg856_out;
SharedReg617_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg617_out;
SharedReg780_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg780_out;
SharedReg428_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg428_out;
SharedReg431_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg431_out;
SharedReg429_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg429_out;
SharedReg830_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg830_out;
SharedReg618_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg618_out;
SharedReg785_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg785_out;
SharedReg832_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg832_out;
SharedReg38_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg38_out;
SharedReg428_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg428_out;
SharedReg66_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg66_out;
SharedReg780_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg780_out;
SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg36_out;
SharedReg834_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg834_out;
SharedReg611_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg611_out;
SharedReg612_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg612_out;
   MUX_Product12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg425_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg423_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg852_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg170_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg765_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg168_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg425_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg42_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg426_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg172_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg174_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg611_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg176_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg44_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg51_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg169_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg426_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg614_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg194_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg855_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg609_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg812_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg613_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg856_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg617_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg423_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg780_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg428_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg431_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg429_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg830_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg618_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg785_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg832_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg38_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg428_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg610_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg66_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg780_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg834_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg611_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg612_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg422_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg36_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product12_0_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product12_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_1_impl_out,
                 X => Delay1No88_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg831_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg831_out;
SharedReg66_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg635_out;
SharedReg742_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg742_out;
SharedReg833_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg833_out;
SharedReg779_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg779_out;
SharedReg474_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg474_out;
SharedReg789_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg789_out;
SharedReg630_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg630_out;
SharedReg835_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg835_out;
SharedReg822_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg822_out;
SharedReg823_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg823_out;
SharedReg824_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg824_out;
SharedReg825_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg825_out;
SharedReg826_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg826_out;
SharedReg827_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg827_out;
SharedReg752_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg760_out;
SharedReg863_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg863_out;
SharedReg715_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg715_out;
SharedReg762_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg762_out;
SharedReg447_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg447_out;
SharedReg718_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg718_out;
SharedReg191_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg191_out;
SharedReg859_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg859_out;
SharedReg766_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg766_out;
SharedReg828_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg828_out;
SharedReg768_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg768_out;
SharedReg814_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg814_out;
SharedReg863_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg863_out;
SharedReg724_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg724_out;
SharedReg725_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg725_out;
SharedReg726_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg726_out;
SharedReg797_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg797_out;
SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg635_out;
SharedReg799_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg799_out;
SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg635_out;
SharedReg801_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg802_out;
SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg635_out;
SharedReg723_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg723_out;
SharedReg630_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg630_out;
SharedReg854_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg854_out;
SharedReg810_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg810_out;
SharedReg753_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg753_out;
SharedReg754_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg758_out;
SharedReg759_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg759_out;
SharedReg723_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg723_out;
SharedReg727_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg727_out;
SharedReg728_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg728_out;
SharedReg729_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg729_out;
SharedReg730_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg730_out;
   MUX_Product12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg831_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg822_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg823_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg824_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg825_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg826_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg827_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg752_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg760_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg863_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg715_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg762_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg447_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg718_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg191_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg859_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg766_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg828_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg768_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg814_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg863_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg742_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg724_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg725_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg726_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg797_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg799_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg801_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg802_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg635_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg833_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg723_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg630_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg854_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg810_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg753_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg754_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg755_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg756_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg757_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg758_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg779_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg759_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg723_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg727_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg728_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg729_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg730_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg474_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg789_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg630_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg835_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product12_1_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_0_out,
                 Y => Delay1No88_out);

SharedReg639_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg639_out;
SharedReg785_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg785_out;
SharedReg832_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg832_out;
SharedReg64_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg64_out;
SharedReg451_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg451_out;
SharedReg92_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg92_out;
SharedReg780_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg780_out;
SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg62_out;
SharedReg834_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg834_out;
SharedReg632_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg632_out;
SharedReg633_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg633_out;
SharedReg448_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg448_out;
SharedReg446_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg446_out;
SharedReg632_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg632_out;
SharedReg630_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg630_out;
SharedReg446_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg446_out;
SharedReg631_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg631_out;
SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg445_out;
SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg445_out;
SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg62_out;
SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg62_out;
SharedReg852_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg852_out;
SharedReg192_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg192_out;
SharedReg765_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg765_out;
SharedReg631_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg631_out;
SharedReg190_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg190_out;
SharedReg448_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg448_out;
SharedReg68_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg68_out;
SharedReg449_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg449_out;
SharedReg468_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg468_out;
SharedReg196_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg196_out;
SharedReg198_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg198_out;
SharedReg70_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg70_out;
SharedReg77_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg77_out;
SharedReg798_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg798_out;
SharedReg635_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg635_out;
SharedReg800_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg800_out;
SharedReg191_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg191_out;
SharedReg449_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg449_out;
SharedReg803_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg803_out;
SharedReg220_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg220_out;
SharedReg772_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg772_out;
SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg445_out;
SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg445_out;
SharedReg213_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg213_out;
SharedReg481_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg481_out;
SharedReg93_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg93_out;
SharedReg91_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg91_out;
SharedReg91_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg91_out;
SharedReg657_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg657_out;
SharedReg656_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg656_out;
SharedReg242_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg242_out;
SharedReg88_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg88_out;
SharedReg210_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg210_out;
SharedReg88_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg88_out;
SharedReg211_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg211_out;
   MUX_Product12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg639_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg785_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg633_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg448_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg446_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg632_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg630_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg446_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg631_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg832_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg852_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg192_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg765_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg631_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg190_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg448_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg68_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg449_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg468_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg64_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg196_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg198_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg70_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg77_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg798_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg635_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg800_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg191_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg449_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg803_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg451_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg220_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg772_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg445_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg213_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg481_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg93_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg91_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg91_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg657_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg92_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg656_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg242_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg88_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg210_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg88_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg211_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg780_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg62_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg834_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg632_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product12_1_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Product12_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_4_impl_out,
                 X => Delay1No90_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg262_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg255_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg255_out;
SharedReg254_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg254_out;
SharedReg257_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg257_out;
SharedReg255_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg255_out;
SharedReg828_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg828_out;
SharedReg718_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg718_out;
SharedReg851_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg851_out;
SharedReg859_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg859_out;
SharedReg776_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
SharedReg717_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg717_out;
SharedReg715_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg715_out;
SharedReg762_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg762_out;
SharedReg741_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg741_out;
SharedReg783_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg783_out;
SharedReg742_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg742_out;
SharedReg727_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg727_out;
SharedReg806_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg806_out;
SharedReg733_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg733_out;
SharedReg782_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg782_out;
SharedReg808_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg808_out;
SharedReg848_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg848_out;
SharedReg818_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg818_out;
SharedReg819_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg819_out;
SharedReg820_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg820_out;
SharedReg827_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg827_out;
SharedReg826_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg826_out;
SharedReg757_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg757_out;
SharedReg824_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg824_out;
SharedReg825_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg825_out;
SharedReg753_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg753_out;
SharedReg756_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg756_out;
SharedReg789_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg789_out;
SharedReg823_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg823_out;
SharedReg822_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg822_out;
SharedReg821_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg821_out;
SharedReg755_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg755_out;
SharedReg754_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg754_out;
SharedReg725_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg725_out;
SharedReg724_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg724_out;
SharedReg771_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg771_out;
SharedReg723_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg723_out;
SharedReg766_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg766_out;
SharedReg863_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg863_out;
   MUX_Product12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_44_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg255_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg717_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg715_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg762_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg741_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg783_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg742_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg727_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg806_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg733_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg782_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg254_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg808_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg848_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg818_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg819_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg820_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg827_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg826_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg757_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg824_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg825_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg257_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg753_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg756_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg789_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg823_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg822_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg821_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg755_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg754_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg725_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg724_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg255_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg771_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg723_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg766_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg863_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_5 => SharedReg828_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg718_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg851_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg859_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product12_4_impl_0_LUT_out,
                 oMux => MUX_Product12_4_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_0_out,
                 Y => Delay1No90_out);

SharedReg258_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg150_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg150_out;
SharedReg258_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg258_out;
SharedReg262_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg144_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg144_out;
SharedReg257_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg257_out;
SharedReg141_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg141_out;
SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg140_out;
SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg140_out;
SharedReg155_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg155_out;
SharedReg260_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg260_out;
SharedReg256_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg256_out;
SharedReg254_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg254_out;
SharedReg264_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg264_out;
SharedReg262_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg262_out;
SharedReg148_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg148_out;
SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg140_out;
SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg514_out;
SharedReg517_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg517_out;
SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg514_out;
SharedReg520_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg520_out;
SharedReg523_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg523_out;
SharedReg704_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg704_out;
SharedReg693_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg693_out;
SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg514_out;
SharedReg702_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg702_out;
SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg698_out;
SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg698_out;
SharedReg515_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg515_out;
SharedReg693_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg693_out;
SharedReg515_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg515_out;
SharedReg695_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg695_out;
SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg698_out;
SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg698_out;
SharedReg696_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg696_out;
SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg694_out;
SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg694_out;
SharedReg517_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg517_out;
SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg694_out;
SharedReg777_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg777_out;
SharedReg775_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg775_out;
SharedReg781_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg781_out;
SharedReg790_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg790_out;
SharedReg765_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg765_out;
   MUX_Product12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_44_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg150_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg260_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg256_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg254_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg264_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg262_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg148_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg517_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg258_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg520_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg523_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg704_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg693_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg514_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg702_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg515_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg693_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg262_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg515_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg695_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg698_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg696_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg517_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg694_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg777_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg144_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg775_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg781_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg790_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg765_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_5 => SharedReg257_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg141_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg140_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg155_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product12_4_impl_1_LUT_out,
                 oMux => MUX_Product12_4_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product22_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_4_impl_out,
                 X => Delay1No92_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast);

SharedReg255_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg255_out;
SharedReg232_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg232_out;
SharedReg118_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg118_out;
SharedReg240_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg240_out;
SharedReg238_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg238_out;
SharedReg499_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg499_out;
SharedReg672_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg672_out;
SharedReg679_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg679_out;
SharedReg677_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg677_out;
SharedReg677_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg677_out;
SharedReg493_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg493_out;
SharedReg520_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg520_out;
SharedReg673_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg673_out;
SharedReg763_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg763_out;
SharedReg805_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg805_out;
SharedReg849_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg849_out;
SharedReg857_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg857_out;
SharedReg861_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg861_out;
SharedReg779_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg779_out;
SharedReg715_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg715_out;
SharedReg762_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg762_out;
SharedReg741_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg741_out;
SharedReg734_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg734_out;
SharedReg742_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg742_out;
SharedReg810_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg810_out;
SharedReg737_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg737_out;
SharedReg807_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg807_out;
SharedReg811_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg811_out;
SharedReg854_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg854_out;
SharedReg847_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg847_out;
SharedReg722_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg722_out;
SharedReg818_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg818_out;
SharedReg819_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg819_out;
SharedReg820_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg820_out;
SharedReg817_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg817_out;
SharedReg827_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg827_out;
SharedReg826_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg826_out;
SharedReg801_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg801_out;
SharedReg824_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg824_out;
SharedReg825_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg825_out;
SharedReg759_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg759_out;
SharedReg802_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg802_out;
SharedReg802_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg802_out;
SharedReg823_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg823_out;
SharedReg836_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg836_out;
SharedReg752_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg752_out;
SharedReg821_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg821_out;
SharedReg799_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg799_out;
SharedReg760_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg760_out;
SharedReg770_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg770_out;
SharedReg771_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg771_out;
SharedReg722_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg722_out;
SharedReg719_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg719_out;
   MUX_Product22_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_53_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg255_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg232_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg493_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg520_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg673_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg763_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg805_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg849_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg857_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg861_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg779_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg715_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg118_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg762_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg741_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg734_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg742_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg810_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg737_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg807_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg811_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg854_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg847_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg240_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg722_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg818_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg819_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg820_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg817_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg827_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg826_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg801_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg824_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg825_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg238_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg759_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg802_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg802_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg823_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg836_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg752_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg821_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg799_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg760_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg770_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg499_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg771_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg722_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg719_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_6 => SharedReg672_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg679_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg677_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg677_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product22_4_impl_0_LUT_out,
                 oMux => MUX_Product22_4_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_0_out,
                 Y => Delay1No92_out);

SharedReg143_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg118_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg118_out;
SharedReg147_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg147_out;
SharedReg235_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg235_out;
SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg114_out;
SharedReg146_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg146_out;
SharedReg242_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg242_out;
SharedReg122_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg122_out;
SharedReg144_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg144_out;
SharedReg494_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg494_out;
SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg673_out;
SharedReg494_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg494_out;
SharedReg501_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg501_out;
SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg491_out;
SharedReg678_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg678_out;
SharedReg497_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg497_out;
SharedReg498_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg498_out;
SharedReg500_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg500_out;
SharedReg676_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg676_out;
SharedReg683_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg683_out;
SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg491_out;
SharedReg681_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg681_out;
SharedReg677_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg677_out;
SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg491_out;
SharedReg495_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg495_out;
SharedReg492_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg492_out;
SharedReg672_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg672_out;
SharedReg699_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg699_out;
SharedReg698_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg698_out;
SharedReg492_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg492_out;
SharedReg674_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg674_out;
SharedReg493_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg493_out;
SharedReg677_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg677_out;
SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg673_out;
SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg673_out;
SharedReg701_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg701_out;
SharedReg497_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg497_out;
SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg673_out;
SharedReg672_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg672_out;
SharedReg772_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg772_out;
SharedReg780_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg780_out;
SharedReg812_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg812_out;
SharedReg856_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg856_out;
SharedReg852_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg852_out;
SharedReg830_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg830_out;
SharedReg796_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg796_out;
SharedReg767_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg767_out;
SharedReg800_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg800_out;
SharedReg790_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg790_out;
SharedReg798_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg798_out;
SharedReg769_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg769_out;
SharedReg766_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg766_out;
   MUX_Product22_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_53_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg494_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg494_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg501_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg678_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg497_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg498_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg500_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg676_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg147_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg683_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg681_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg677_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg491_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg495_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg492_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg672_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg699_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg698_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg235_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg492_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg674_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg493_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg677_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg701_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg497_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg673_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg672_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg772_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg780_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg812_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg856_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg852_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg830_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg796_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg767_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg800_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg790_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg114_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg798_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg769_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg766_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_6 => SharedReg146_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg242_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg122_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg144_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product22_4_impl_1_LUT_out,
                 oMux => MUX_Product22_4_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product6_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_0_impl_out,
                 X => Delay1No94_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg425_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg425_out;
SharedReg838_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg838_out;
SharedReg611_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg611_out;
SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg609_out;
SharedReg841_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg841_out;
SharedReg610_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg610_out;
SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg609_out;
SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg609_out;
SharedReg36_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg36_out;
SharedReg716_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg716_out;
SharedReg717_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg717_out;
SharedReg805_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg805_out;
SharedReg719_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg719_out;
SharedReg861_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg861_out;
SharedReg172_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg172_out;
SharedReg40_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg40_out;
SharedReg722_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg722_out;
SharedReg815_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg815_out;
SharedReg723_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg723_out;
SharedReg174_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg174_out;
SharedReg770_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg770_out;
SharedReg771_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg771_out;
SharedReg797_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg797_out;
SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg614_out;
SharedReg799_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg799_out;
SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg614_out;
SharedReg801_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg802_out;
SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg614_out;
SharedReg723_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg723_out;
SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg609_out;
SharedReg854_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg854_out;
SharedReg810_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg810_out;
SharedReg753_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg753_out;
SharedReg754_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg754_out;
SharedReg755_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg755_out;
SharedReg756_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg756_out;
SharedReg757_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg757_out;
SharedReg758_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg758_out;
SharedReg759_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg759_out;
SharedReg843_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg843_out;
SharedReg727_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg727_out;
SharedReg728_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg728_out;
SharedReg729_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg729_out;
SharedReg730_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg730_out;
SharedReg731_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg731_out;
SharedReg732_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg732_out;
SharedReg808_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg808_out;
SharedReg635_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg635_out;
SharedReg734_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg734_out;
SharedReg850_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg850_out;
SharedReg843_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg843_out;
SharedReg194_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg194_out;
SharedReg738_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg738_out;
SharedReg739_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg739_out;
SharedReg740_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg740_out;
   MUX_Product6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg425_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg838_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg717_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg805_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg719_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg861_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg172_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg40_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg722_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg815_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg723_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg174_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg611_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg770_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg771_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg797_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg799_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg801_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg802_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg614_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg723_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg854_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg810_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg753_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg754_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg755_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg756_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg757_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg758_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg759_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg841_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg843_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg727_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg728_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg729_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg730_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg731_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg732_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg808_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg635_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg734_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg610_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg850_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg843_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg194_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg738_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg739_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg740_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg609_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg36_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg716_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product6_0_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_0_out,
                 Y => Delay1No94_out);

SharedReg837_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg837_out;
SharedReg423_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg423_out;
SharedReg839_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg839_out;
SharedReg840_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg840_out;
SharedReg423_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg796_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg796_out;
SharedReg760_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg760_out;
SharedReg863_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg863_out;
SharedReg761_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg761_out;
SharedReg166_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg166_out;
SharedReg37_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg37_out;
SharedReg424_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg424_out;
SharedReg615_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg615_out;
SharedReg610_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg610_out;
SharedReg766_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg766_out;
SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg767_out;
SharedReg432_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg432_out;
SharedReg429_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg429_out;
SharedReg176_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg176_out;
SharedReg769_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg769_out;
SharedReg176_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg176_out;
SharedReg44_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg44_out;
SharedReg51_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg51_out;
SharedReg798_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg798_out;
SharedReg614_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg614_out;
SharedReg800_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg800_out;
SharedReg169_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg169_out;
SharedReg426_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg426_out;
SharedReg803_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg803_out;
SharedReg198_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg198_out;
SharedReg772_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg772_out;
SharedReg422_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg422_out;
SharedReg191_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg191_out;
SharedReg458_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg458_out;
SharedReg67_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg67_out;
SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg65_out;
SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg65_out;
SharedReg636_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg636_out;
SharedReg66_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg66_out;
SharedReg658_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg658_out;
SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg62_out;
SharedReg188_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg188_out;
SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg62_out;
SharedReg189_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg189_out;
SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg62_out;
SharedReg189_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg189_out;
SharedReg634_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg634_out;
SharedReg813_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg813_out;
SharedReg69_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg69_out;
SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg638_out;
SharedReg679_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg679_out;
SharedReg781_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg781_out;
SharedReg195_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg195_out;
SharedReg72_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg72_out;
SharedReg196_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg196_out;
   MUX_Product6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg837_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg423_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg37_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg424_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg615_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg610_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg766_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg767_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg432_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg429_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg176_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg769_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg839_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg176_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg44_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg51_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg798_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg614_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg800_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg169_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg426_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg803_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg198_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg840_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg772_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg422_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg422_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg191_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg458_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg67_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg65_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg636_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg66_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg423_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg658_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg188_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg189_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg189_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg634_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg813_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg69_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg796_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg679_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg781_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg195_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg72_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg196_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg760_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg863_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg761_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg166_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Product6_0_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product6_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_4_impl_out,
                 X => Delay1No96_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg144_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg144_out;
SharedReg140_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg140_out;
SharedReg144_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg144_out;
SharedReg262_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg260_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg260_out;
SharedReg517_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg517_out;
SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg693_out;
SharedReg522_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg522_out;
SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg693_out;
SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg693_out;
SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg698_out;
SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg698_out;
SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg693_out;
SharedReg695_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg695_out;
SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg698_out;
SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg693_out;
SharedReg694_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg694_out;
SharedReg805_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg805_out;
SharedReg849_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg849_out;
SharedReg857_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg857_out;
SharedReg861_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg861_out;
SharedReg742_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg742_out;
SharedReg810_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg810_out;
SharedReg737_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg737_out;
SharedReg807_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg807_out;
SharedReg811_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg811_out;
SharedReg854_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg854_out;
SharedReg831_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg831_out;
SharedReg817_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg817_out;
SharedReg833_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg833_out;
SharedReg841_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg841_out;
SharedReg801_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg801_out;
SharedReg838_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg838_out;
SharedReg797_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg797_out;
SharedReg789_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg789_out;
SharedReg835_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg835_out;
SharedReg799_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg799_out;
SharedReg770_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg770_out;
SharedReg716_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg716_out;
SharedReg723_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg723_out;
SharedReg719_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg719_out;
   MUX_Product6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_41_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg144_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg140_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg695_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg698_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg694_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg805_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg849_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg857_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg144_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg861_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg742_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg810_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg737_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg807_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg811_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg854_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg831_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg817_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg833_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg262_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg841_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg801_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg838_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg797_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg789_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg835_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg799_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg770_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg716_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg723_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg260_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg719_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_5 => SharedReg517_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg522_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg693_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product6_4_impl_0_LUT_out,
                 oMux => MUX_Product6_4_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_0_out,
                 Y => Delay1No96_out);

SharedReg142_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg257_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg257_out;
SharedReg155_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg155_out;
SharedReg140_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg140_out;
SharedReg264_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg264_out;
SharedReg254_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg254_out;
SharedReg264_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg264_out;
SharedReg699_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg699_out;
SharedReg520_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg520_out;
SharedReg521_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg521_out;
SharedReg523_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg523_out;
SharedReg697_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg697_out;
SharedReg514_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg514_out;
SharedReg702_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg702_out;
SharedReg514_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg514_out;
SharedReg515_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg515_out;
SharedReg515_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg515_out;
SharedReg516_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg516_out;
SharedReg698_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg698_out;
SharedReg695_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg695_out;
SharedReg694_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg694_out;
SharedReg520_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg520_out;
SharedReg694_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_23_cast <= SharedReg694_out;
SharedReg693_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg693_out;
SharedReg855_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg855_out;
SharedReg761_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg761_out;
SharedReg785_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg785_out;
SharedReg772_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg772_out;
SharedReg812_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg812_out;
SharedReg832_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg832_out;
SharedReg830_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg830_out;
SharedReg840_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg840_out;
SharedReg839_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg839_out;
SharedReg767_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg767_out;
SharedReg800_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg800_out;
SharedReg837_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg837_out;
SharedReg834_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg834_out;
SharedReg798_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg798_out;
SharedReg769_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg769_out;
SharedReg766_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg766_out;
SharedReg863_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg863_out;
   MUX_Product6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_41_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg523_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg697_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg514_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg702_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg514_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg515_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg515_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg516_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg698_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg695_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg155_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg694_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg520_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg694_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg693_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg855_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg761_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg785_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg772_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg812_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg832_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg140_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg830_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg840_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg839_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg767_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg800_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg837_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg834_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg798_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg769_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg766_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg264_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg863_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_5 => SharedReg254_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg264_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg699_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg520_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg521_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product6_4_impl_1_LUT_out,
                 oMux => MUX_Product6_4_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Subtract9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_0_impl_out,
                 X => Delay1No98_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg623_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg623_out;
SharedReg1_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg13_out;
SharedReg543_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg543_out;
SharedReg283_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg283_out;
SharedReg276_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg276_out;
SharedReg544_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg544_out;
SharedReg47_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg47_out;
SharedReg433_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg433_out;
SharedReg52_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg52_out;
SharedReg624_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg624_out;
SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg537_out;
SharedReg182_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg182_out;
SharedReg59_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg59_out;
SharedReg586_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg586_out;
SharedReg628_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg628_out;
SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg537_out;
SharedReg186_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg186_out;
SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg537_out;
SharedReg170_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg170_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg166_out;
SharedReg177_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg177_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg166_out;
SharedReg429_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg429_out;
SharedReg176_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg176_out;
SharedReg432_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg432_out;
SharedReg616_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg616_out;
SharedReg282_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg282_out;
SharedReg543_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg543_out;
SharedReg541_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg541_out;
SharedReg281_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg281_out;
SharedReg50_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg50_out;
SharedReg422_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg422_out;
SharedReg37_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg37_out;
SharedReg611_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg611_out;
SharedReg169_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg169_out;
SharedReg544_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg544_out;
SharedReg40_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg40_out;
SharedReg171_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg171_out;
SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg537_out;
SharedReg428_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg428_out;
SharedReg423_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg423_out;
SharedReg39_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg39_out;
SharedReg45_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg45_out;
SharedReg278_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg278_out;
SharedReg172_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg172_out;
SharedReg361_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg361_out;
SharedReg358_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg358_out;
SharedReg176_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg176_out;
SharedReg37_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg37_out;
   MUX_Subtract9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg623_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg283_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg276_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg544_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg47_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg433_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg52_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg624_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg182_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg59_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg3_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg586_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg628_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg186_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg170_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg166_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg177_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg166_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg429_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg17_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg176_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg432_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg616_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg282_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg543_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg541_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg281_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg50_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg422_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg37_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg6_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg611_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg169_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg544_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg40_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg171_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg537_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg428_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg423_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg39_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg45_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg11_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg278_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg172_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg361_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg358_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg176_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg37_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg12_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg13_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg543_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_0_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_0_out,
                 Y => Delay1No98_out);

SharedReg443_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg443_out;
SharedReg19_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg31_out;
SharedReg545_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg545_out;
SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg591_out;
SharedReg586_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg586_out;
SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg591_out;
SharedReg178_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg178_out;
SharedReg621_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg621_out;
SharedReg176_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg176_out;
SharedReg622_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg622_out;
SharedReg363_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg363_out;
SharedReg180_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg180_out;
SharedReg61_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg61_out;
SharedReg594_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg594_out;
SharedReg629_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg629_out;
SharedReg589_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg589_out;
SharedReg187_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg187_out;
SharedReg587_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg587_out;
SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg167_out;
SharedReg170_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg170_out;
SharedReg36_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg36_out;
SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg167_out;
SharedReg609_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg609_out;
SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg167_out;
SharedReg423_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg423_out;
SharedReg429_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg429_out;
Delay25No35_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_34_cast <= Delay25No35_out;
SharedReg592_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg592_out;
SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg591_out;
SharedReg589_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg589_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg166_out;
SharedReg437_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg437_out;
SharedReg55_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg55_out;
SharedReg626_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg626_out;
SharedReg183_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg183_out;
SharedReg537_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg537_out;
SharedReg56_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg56_out;
SharedReg184_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg184_out;
SharedReg538_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg538_out;
SharedReg440_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg440_out;
SharedReg609_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg609_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg166_out;
SharedReg57_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg57_out;
SharedReg537_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg537_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg166_out;
SharedReg538_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg538_out;
SharedReg542_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg542_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg166_out;
SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg166_out;
   MUX_Subtract9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg443_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg586_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg178_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg621_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg176_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg622_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg363_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg180_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg61_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg594_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg629_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg589_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg187_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg587_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg170_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg36_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg609_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg35_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg167_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg423_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg429_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => Delay25No35_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg592_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg591_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg589_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg437_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg55_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg626_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg183_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg537_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg56_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg184_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg538_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg440_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg609_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg57_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg29_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg537_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg538_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg542_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg166_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg30_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg34_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg31_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg545_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_0_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Subtract9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_1_impl_out,
                 X => Delay1No100_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg370_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg370_out;
SharedReg451_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg451_out;
SharedReg446_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg446_out;
SharedReg65_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg65_out;
SharedReg71_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg71_out;
SharedReg588_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg588_out;
SharedReg194_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg194_out;
SharedReg373_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg373_out;
SharedReg370_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg370_out;
SharedReg198_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg198_out;
SharedReg63_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg63_out;
SharedReg644_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg644_out;
SharedReg1_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg13_out;
SharedReg555_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg555_out;
SharedReg294_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg294_out;
SharedReg287_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg287_out;
SharedReg556_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg556_out;
SharedReg73_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg73_out;
SharedReg456_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg456_out;
SharedReg78_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg78_out;
SharedReg645_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg645_out;
SharedReg550_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg550_out;
SharedReg204_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg204_out;
SharedReg85_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg85_out;
SharedReg322_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg322_out;
SharedReg649_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg649_out;
SharedReg537_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg537_out;
SharedReg208_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg208_out;
SharedReg550_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg550_out;
SharedReg192_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg192_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg188_out;
SharedReg199_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg199_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg188_out;
SharedReg452_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg452_out;
SharedReg198_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg198_out;
SharedReg455_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg455_out;
SharedReg637_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg637_out;
SharedReg591_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg591_out;
SharedReg376_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg376_out;
SharedReg374_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg374_out;
SharedReg590_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg590_out;
SharedReg76_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg76_out;
SharedReg445_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg445_out;
SharedReg63_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg63_out;
SharedReg632_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg632_out;
SharedReg191_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg191_out;
SharedReg377_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg377_out;
SharedReg66_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg66_out;
SharedReg193_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg193_out;
   MUX_Subtract9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg370_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg451_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg63_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg644_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg3_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg17_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg6_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg11_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg12_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg16_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg13_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg446_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg555_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg294_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg287_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg556_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg73_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg456_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg78_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg645_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg550_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg204_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg65_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg85_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg322_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg649_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg537_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg208_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg550_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg192_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg188_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg199_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg188_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg71_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg452_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg198_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg455_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg637_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg591_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg376_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg374_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg590_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg76_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg445_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg588_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg63_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg632_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg191_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg377_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg66_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg193_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg194_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg373_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg370_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg198_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_1_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_0_out,
                 Y => Delay1No100_out);

SharedReg538_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg538_out;
SharedReg463_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg463_out;
SharedReg630_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg630_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg188_out;
SharedReg83_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg83_out;
SharedReg550_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg550_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg188_out;
SharedReg551_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg551_out;
SharedReg375_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg375_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg188_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg188_out;
SharedReg466_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg466_out;
SharedReg19_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_17_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg31_out;
SharedReg557_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg557_out;
SharedReg327_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg327_out;
SharedReg322_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg322_out;
SharedReg327_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg327_out;
SharedReg200_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg200_out;
SharedReg642_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg642_out;
SharedReg198_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg198_out;
SharedReg643_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg643_out;
SharedReg375_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg375_out;
SharedReg202_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg202_out;
SharedReg87_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg87_out;
SharedReg330_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg330_out;
SharedReg650_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg650_out;
SharedReg325_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg325_out;
SharedReg209_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg209_out;
SharedReg323_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg323_out;
SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg189_out;
SharedReg192_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg192_out;
SharedReg62_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg62_out;
SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg189_out;
SharedReg630_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg630_out;
SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg189_out;
SharedReg446_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg446_out;
SharedReg452_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg452_out;
Delay25No36_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_45_cast <= Delay25No36_out;
SharedReg556_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg556_out;
SharedReg555_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg555_out;
SharedReg553_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg553_out;
SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg188_out;
SharedReg460_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg460_out;
SharedReg81_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg81_out;
SharedReg647_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg647_out;
SharedReg205_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg205_out;
SharedReg370_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg370_out;
SharedReg82_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg82_out;
SharedReg206_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg206_out;
   MUX_Subtract9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg538_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg463_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg466_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg21_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg35_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg24_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg29_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg30_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg34_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg31_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg630_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg557_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg327_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg322_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg327_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg200_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg642_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg198_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg643_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg375_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg202_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg87_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg330_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg650_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg325_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg209_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg323_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg192_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg62_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg83_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg630_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg189_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg446_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg452_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => Delay25No36_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg556_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg555_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg553_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg460_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg550_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg81_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg647_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg205_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg370_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg82_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg206_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg551_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg375_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg188_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_1_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Subtract9_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_2_impl_out,
                 X => Delay1No102_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg304_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg302_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg302_out;
SharedReg554_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg554_out;
SharedReg102_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg102_out;
SharedReg468_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg468_out;
SharedReg89_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg89_out;
SharedReg653_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg653_out;
SharedReg213_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg213_out;
SharedReg305_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg305_out;
SharedReg92_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg92_out;
SharedReg215_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg215_out;
SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg383_out;
SharedReg474_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg474_out;
SharedReg469_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg469_out;
SharedReg91_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg91_out;
SharedReg97_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg97_out;
SharedReg324_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg324_out;
SharedReg216_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg216_out;
SharedReg386_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg386_out;
SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg383_out;
SharedReg220_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg220_out;
SharedReg89_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg89_out;
SharedReg665_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg665_out;
SharedReg1_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg13_out;
SharedReg338_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg338_out;
SharedReg305_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg305_out;
SharedReg287_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg287_out;
SharedReg339_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg339_out;
SharedReg99_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg99_out;
SharedReg479_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg479_out;
SharedReg104_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg104_out;
SharedReg666_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg666_out;
SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg383_out;
SharedReg226_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg226_out;
SharedReg111_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg111_out;
SharedReg333_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg333_out;
SharedReg670_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg670_out;
SharedReg370_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg370_out;
SharedReg230_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg230_out;
SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg383_out;
SharedReg214_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg214_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg210_out;
SharedReg221_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg221_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg210_out;
SharedReg475_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg475_out;
SharedReg220_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg220_out;
SharedReg478_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg478_out;
SharedReg658_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg658_out;
SharedReg555_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg555_out;
   MUX_Subtract9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg302_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg215_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg474_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg469_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg91_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg97_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg324_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg216_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg386_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg554_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg220_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg89_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg665_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg1_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg3_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg17_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg6_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg11_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg12_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg16_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg102_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg13_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg338_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg305_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg287_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg339_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg99_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg479_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg104_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg666_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg468_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg226_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg111_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg333_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg670_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg370_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg230_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg383_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg214_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg210_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg221_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg89_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg210_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg475_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg220_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg478_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg658_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg555_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg653_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg213_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg305_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg92_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_2_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_2_impl_0_out,
                 Y => Delay1No102_out);

SharedReg390_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg389_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg325_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg325_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg210_out;
SharedReg483_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg483_out;
SharedReg107_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg107_out;
SharedReg668_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg668_out;
SharedReg227_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg227_out;
SharedReg383_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg383_out;
SharedReg108_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg108_out;
SharedReg228_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg228_out;
SharedReg551_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg486_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg486_out;
SharedReg651_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg651_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg210_out;
SharedReg109_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg109_out;
SharedReg333_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg333_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg210_out;
SharedReg334_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg334_out;
SharedReg388_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg388_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg210_out;
SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg210_out;
SharedReg489_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg489_out;
SharedReg19_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg31_out;
SharedReg340_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg340_out;
SharedReg316_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg316_out;
SharedReg322_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg322_out;
SharedReg316_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg316_out;
SharedReg222_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg222_out;
SharedReg663_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg663_out;
SharedReg220_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg220_out;
SharedReg664_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg664_out;
SharedReg388_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg388_out;
SharedReg224_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg224_out;
SharedReg113_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg113_out;
SharedReg318_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg318_out;
SharedReg671_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg671_out;
SharedReg336_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg336_out;
SharedReg231_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg231_out;
SharedReg334_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg334_out;
SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg211_out;
SharedReg214_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg214_out;
SharedReg88_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg88_out;
SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg211_out;
SharedReg651_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg651_out;
SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg211_out;
SharedReg469_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg469_out;
SharedReg475_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg475_out;
SharedReg321_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg321_out;
   MUX_Subtract9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg228_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg486_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg651_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg109_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg333_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg334_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg388_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg325_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg489_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg19_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg21_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg35_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg24_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg29_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg30_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg34_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg210_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg31_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg340_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg316_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg322_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg316_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg222_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg663_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg220_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg664_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg388_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg483_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg224_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg113_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg318_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg671_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg336_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg231_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg334_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg214_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg88_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg107_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg651_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg211_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg469_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg475_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg321_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg668_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg227_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg383_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg108_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_2_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_2_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Subtract9_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_3_impl_out,
                 X => Delay1No104_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast);

SharedReg252_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg252_out;
SharedReg396_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg236_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg243_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg243_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg232_out;
SharedReg498_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg498_out;
SharedReg242_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg242_out;
SharedReg501_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg501_out;
SharedReg679_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg679_out;
SharedReg338_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg338_out;
SharedReg402_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg402_out;
SharedReg400_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg400_out;
SharedReg337_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg337_out;
SharedReg128_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg128_out;
SharedReg491_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg491_out;
SharedReg115_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg115_out;
SharedReg674_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg674_out;
SharedReg235_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg235_out;
SharedReg403_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg403_out;
SharedReg118_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg118_out;
SharedReg237_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg237_out;
SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg574_out;
SharedReg497_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg497_out;
SharedReg492_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg492_out;
SharedReg117_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg117_out;
SharedReg123_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg123_out;
SharedReg312_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg312_out;
SharedReg238_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg238_out;
SharedReg577_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg577_out;
SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg574_out;
SharedReg242_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg242_out;
SharedReg115_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg115_out;
SharedReg686_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg686_out;
SharedReg1_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg13_out;
SharedReg351_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg351_out;
SharedReg403_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg403_out;
SharedReg322_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg322_out;
SharedReg581_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg581_out;
SharedReg125_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg125_out;
SharedReg502_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg502_out;
SharedReg130_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg130_out;
SharedReg687_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg687_out;
SharedReg396_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg396_out;
SharedReg248_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg248_out;
SharedReg137_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg137_out;
SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg574_out;
SharedReg691_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg691_out;
SharedReg370_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg370_out;
   MUX_Subtract9_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg252_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg338_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg402_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg400_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg337_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg128_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg491_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg115_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg674_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg235_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg403_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg236_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg118_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg237_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg497_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg492_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg117_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg123_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg312_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg238_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg577_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg232_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg242_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg115_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg686_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg1_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg3_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg17_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg6_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg11_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg12_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg243_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg16_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg13_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg351_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg403_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg322_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg581_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg125_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg502_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg130_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg687_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg232_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg396_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg248_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg137_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg574_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg691_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg370_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg498_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg242_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg501_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg679_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_3_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_3_impl_0_out,
                 Y => Delay1No104_out);

SharedReg253_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg253_out;
SharedReg575_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg575_out;
SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg233_out;
SharedReg236_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg236_out;
SharedReg114_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg114_out;
SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg233_out;
SharedReg672_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg672_out;
SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg233_out;
SharedReg492_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg492_out;
SharedReg498_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg498_out;
SharedReg357_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg357_out;
SharedReg581_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg581_out;
SharedReg580_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg580_out;
SharedReg314_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg314_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg232_out;
SharedReg506_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg506_out;
SharedReg133_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg133_out;
SharedReg689_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_18_cast <= SharedReg689_out;
SharedReg249_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg249_out;
SharedReg574_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg574_out;
SharedReg134_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg134_out;
SharedReg250_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg250_out;
SharedReg334_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_23_cast <= SharedReg334_out;
SharedReg509_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg509_out;
SharedReg672_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg672_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg232_out;
SharedReg135_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg135_out;
SharedReg345_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg345_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg232_out;
SharedReg346_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg346_out;
SharedReg579_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg579_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg232_out;
SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg232_out;
SharedReg512_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg512_out;
SharedReg19_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg31_out;
SharedReg353_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg353_out;
SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg351_out;
SharedReg333_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg333_out;
SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_46_cast <= SharedReg351_out;
SharedReg244_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg244_out;
SharedReg684_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg684_out;
SharedReg242_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg242_out;
SharedReg685_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg685_out;
SharedReg401_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg401_out;
SharedReg246_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg246_out;
SharedReg139_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg139_out;
SharedReg354_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg354_out;
SharedReg692_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg692_out;
SharedReg578_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg578_out;
   MUX_Subtract9_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg253_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg575_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg357_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg581_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg580_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg314_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg506_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg133_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg689_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg249_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg574_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg134_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg250_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg334_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg509_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg672_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg135_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg345_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg346_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg236_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg579_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg232_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg512_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg19_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg21_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg35_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg24_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg29_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg30_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg114_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg34_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg31_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg353_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg333_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg351_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg244_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg684_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg242_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg685_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg401_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg246_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg139_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg354_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg692_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg578_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg672_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg233_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg492_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg498_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_3_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_3_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Subtract9_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_4_impl_out,
                 X => Delay1No106_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast);

SharedReg345_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg345_out;
SharedReg570_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg570_out;
SharedReg151_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg525_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg525_out;
SharedReg156_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg156_out;
SharedReg708_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg708_out;
SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg563_out;
SharedReg270_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg270_out;
SharedReg163_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg163_out;
SharedReg410_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg410_out;
SharedReg712_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg712_out;
SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg563_out;
SharedReg274_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg274_out;
SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg563_out;
SharedReg258_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_15_cast <= SharedReg258_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_16_cast <= SharedReg254_out;
SharedReg265_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_17_cast <= SharedReg265_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_18_cast <= SharedReg254_out;
SharedReg521_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_19_cast <= SharedReg521_out;
SharedReg264_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_20_cast <= SharedReg264_out;
SharedReg524_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_21_cast <= SharedReg524_out;
SharedReg700_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_22_cast <= SharedReg700_out;
SharedReg351_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_23_cast <= SharedReg351_out;
SharedReg569_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_24_cast <= SharedReg569_out;
SharedReg349_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_25_cast <= SharedReg349_out;
SharedReg401_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_26_cast <= SharedReg401_out;
SharedReg154_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_27_cast <= SharedReg154_out;
SharedReg514_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_28_cast <= SharedReg514_out;
SharedReg141_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_29_cast <= SharedReg141_out;
SharedReg695_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_30_cast <= SharedReg695_out;
SharedReg257_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_31_cast <= SharedReg257_out;
SharedReg570_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_32_cast <= SharedReg570_out;
SharedReg144_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_33_cast <= SharedReg144_out;
SharedReg259_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_34_cast <= SharedReg259_out;
SharedReg598_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_35_cast <= SharedReg598_out;
SharedReg520_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_36_cast <= SharedReg520_out;
SharedReg515_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_37_cast <= SharedReg515_out;
SharedReg143_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_38_cast <= SharedReg143_out;
SharedReg149_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_39_cast <= SharedReg149_out;
SharedReg412_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_40_cast <= SharedReg412_out;
SharedReg260_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_41_cast <= SharedReg260_out;
SharedReg566_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_42_cast <= SharedReg566_out;
SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_43_cast <= SharedReg563_out;
SharedReg264_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_44_cast <= SharedReg264_out;
SharedReg141_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_45_cast <= SharedReg141_out;
SharedReg707_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_46_cast <= SharedReg707_out;
SharedReg1_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_47_cast <= SharedReg1_out;
SharedReg3_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_48_cast <= SharedReg3_out;
SharedReg17_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_49_cast <= SharedReg17_out;
SharedReg6_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_50_cast <= SharedReg6_out;
SharedReg11_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_51_cast <= SharedReg11_out;
SharedReg12_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_52_cast <= SharedReg12_out;
SharedReg16_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_53_cast <= SharedReg16_out;
SharedReg13_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_54_cast <= SharedReg13_out;
SharedReg569_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_55_cast <= SharedReg569_out;
SharedReg352_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_56_cast <= SharedReg352_out;
   MUX_Subtract9_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg345_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg570_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg712_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg274_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg258_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg254_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg265_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg254_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg521_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg264_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg151_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg524_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg700_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg351_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg569_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg349_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg401_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg154_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg514_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg141_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg695_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg525_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg257_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg570_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg144_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg259_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg598_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg520_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg515_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg143_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg149_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg412_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg156_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg260_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg566_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg264_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg141_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg707_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg1_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg3_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg17_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg6_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg708_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg11_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg12_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg16_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg13_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg569_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg352_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg563_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg270_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg163_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg410_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_4_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_4_impl_0_out,
                 Y => Delay1No106_out);

SharedReg598_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg598_out;
SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg604_out;
SharedReg266_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg266_out;
SharedReg705_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg705_out;
SharedReg264_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg264_out;
SharedReg706_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg706_out;
SharedReg414_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg414_out;
SharedReg268_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg268_out;
SharedReg165_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg165_out;
SharedReg342_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg342_out;
SharedReg713_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg713_out;
SharedReg602_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg602_out;
SharedReg275_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg275_out;
SharedReg599_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg599_out;
SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_15_cast <= SharedReg255_out;
SharedReg258_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_16_cast <= SharedReg258_out;
SharedReg140_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_17_cast <= SharedReg140_out;
SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_18_cast <= SharedReg255_out;
SharedReg693_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_19_cast <= SharedReg693_out;
SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_20_cast <= SharedReg255_out;
SharedReg515_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_21_cast <= SharedReg515_out;
SharedReg521_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_22_cast <= SharedReg521_out;
Delay25No39_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_23_cast <= Delay25No39_out;
SharedReg605_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_24_cast <= SharedReg605_out;
SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_25_cast <= SharedReg604_out;
SharedReg349_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_26_cast <= SharedReg349_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_27_cast <= SharedReg254_out;
SharedReg529_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_28_cast <= SharedReg529_out;
SharedReg159_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_29_cast <= SharedReg159_out;
SharedReg710_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_30_cast <= SharedReg710_out;
SharedReg271_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_31_cast <= SharedReg271_out;
SharedReg410_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_32_cast <= SharedReg410_out;
SharedReg160_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_33_cast <= SharedReg160_out;
SharedReg272_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_34_cast <= SharedReg272_out;
SharedReg575_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_35_cast <= SharedReg575_out;
SharedReg532_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_36_cast <= SharedReg532_out;
SharedReg693_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_37_cast <= SharedReg693_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_38_cast <= SharedReg254_out;
SharedReg161_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_39_cast <= SharedReg161_out;
SharedReg598_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_40_cast <= SharedReg598_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_41_cast <= SharedReg254_out;
SharedReg599_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_42_cast <= SharedReg599_out;
SharedReg603_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_43_cast <= SharedReg603_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_44_cast <= SharedReg254_out;
SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_45_cast <= SharedReg254_out;
SharedReg535_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_46_cast <= SharedReg535_out;
SharedReg19_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_47_cast <= SharedReg19_out;
SharedReg21_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_48_cast <= SharedReg21_out;
SharedReg35_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_49_cast <= SharedReg35_out;
SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_50_cast <= SharedReg24_out;
SharedReg29_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_51_cast <= SharedReg29_out;
SharedReg30_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_52_cast <= SharedReg30_out;
SharedReg34_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_53_cast <= SharedReg34_out;
SharedReg31_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_54_cast <= SharedReg31_out;
SharedReg606_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_55_cast <= SharedReg606_out;
SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_56_cast <= SharedReg604_out;
   MUX_Subtract9_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_56_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg598_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg713_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg602_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg275_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg599_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg258_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg140_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg693_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg255_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg266_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg515_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg521_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay25No39_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg605_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg349_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg529_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg159_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg710_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg705_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg271_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg410_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg160_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg272_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg575_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg532_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg693_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg161_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg598_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg264_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg599_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg603_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg254_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg535_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg19_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg21_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg35_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg706_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg29_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg30_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg34_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg31_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg606_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg604_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_56_cast,
                 iS_6 => SharedReg414_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg268_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg165_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg342_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount561_out,
                 oMux => MUX_Subtract9_4_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_4_impl_1_out,
                 Y => Delay1No107_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay19No14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => Delay19No14_out);

   Delay19No19_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => Delay19No19_out);

   Delay61No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay61No_out);

   Delay61No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => Delay61No1_out);

   Delay61No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => Delay61No2_out);

   Delay61No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => Delay61No3_out);

   Delay61No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay61No4_out);

   Delay61No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => Delay61No5_out);

   Delay61No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => Delay61No6_out);

   Delay61No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => Delay61No7_out);

   Delay61No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => Delay61No8_out);

   Delay61No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => Delay61No9_out);

   Delay25No15_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => Delay25No15_out);

   Delay25No16_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => Delay25No16_out);

   Delay25No17_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => Delay25No17_out);

   Delay25No20_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => Delay25No20_out);

   Delay25No21_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => Delay25No21_out);

   Delay25No22_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => Delay25No22_out);

   Delay25No30_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => Delay25No30_out);

   Delay25No31_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => Delay25No31_out);

   Delay25No32_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => Delay25No32_out);

   Delay25No35_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => Delay25No35_out);

   Delay25No36_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => Delay25No36_out);

   Delay25No39_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => Delay25No39_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Product4_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product4_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product4_3_impl_0_LUT_out);

   MUX_Product4_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product4_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product4_3_impl_1_LUT_out);

   MUX_Product11_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product11_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product11_4_impl_0_LUT_out);

   MUX_Product11_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product11_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product11_4_impl_1_LUT_out);

   MUX_Product21_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product21_3_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product21_3_impl_0_LUT_out);

   MUX_Product21_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product21_3_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product21_3_impl_1_LUT_out);

   MUX_Product31_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product31_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product31_4_impl_0_LUT_out);

   MUX_Product31_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product31_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product31_4_impl_1_LUT_out);

   MUX_Product12_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product12_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product12_4_impl_0_LUT_out);

   MUX_Product12_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product12_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product12_4_impl_1_LUT_out);

   MUX_Product22_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product22_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product22_4_impl_0_LUT_out);

   MUX_Product22_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product22_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product22_4_impl_1_LUT_out);

   MUX_Product6_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product6_4_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product6_4_impl_0_LUT_out);

   MUX_Product6_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product6_4_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount561_out,
                 Output => MUX_Product6_4_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_3_impl_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_4_impl_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_1_impl_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_2_impl_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_3_impl_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_4_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_0_impl_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_1_impl_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_4_impl_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_4_impl_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_0_impl_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_4_impl_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_0_impl_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_1_impl_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_2_impl_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_3_impl_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_4_impl_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg863_out);
end architecture;

