--------------------------------------------------------------------------------
--                         ModuloCounter_6_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_6_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of ModuloCounter_6_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(2 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 5 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1463306_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1463308)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1463306_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1463306_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1463311
--                  (IntAdderAlternative_27_f250_uid1463315)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1463311 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1463311 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1463318
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1463318 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1463318 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1463321
--                   (IntAdderClassical_34_f250_uid1463323)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1463321 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1463321 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1463306
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1463306 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1463306 is
   component FPAdd_8_23_uid1463306_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1463311 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1463318 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1463321 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1463306_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1463311  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1463318  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1463321  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid1463306 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid1463306  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_6_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_6_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_6_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1466079
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1466079 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1466079 is
signal XX_m1466080 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m1466080 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m1466080 <= X ;
   YY_m1466080 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid1466083
--                   (IntAdderClassical_33_f500_uid1466085)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid1466083 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid1466083 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1466079 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid1466083 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid1466079  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid1466083  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid1466408_RightShifter
--                (RightShifter_24_by_max_26_F250_uid1466410)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1466408_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1466408_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid1466413
--                  (IntAdderAlternative_27_f250_uid1466417)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid1466413 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid1466413 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid1466420
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid1466420 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid1466420 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid1466423
--                   (IntAdderClassical_34_f250_uid1466425)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid1466423 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid1466423 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid1466408
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid1466408 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid1466408 is
   component FPAdd_8_23_uid1466408_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid1466413 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid1466420 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid1466423 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid1466408_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid1466413  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid1466420  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid1466423  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid1466408 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid1466408  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "010" when "000",
      "011" when "001",
      "000" when "010",
      "100" when "011",
      "000" when "100",
      "001" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "010" when "000",
      "011" when "001",
      "000" when "010",
      "100" when "011",
      "000" when "100",
      "001" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "010" when "000",
      "011" when "001",
      "000" when "010",
      "100" when "011",
      "000" when "100",
      "001" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "010" when "000",
      "011" when "001",
      "000" when "010",
      "100" when "011",
      "000" when "100",
      "001" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "010" when "000",
      "011" when "001",
      "000" when "010",
      "100" when "011",
      "000" when "100",
      "001" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "001" when "000",
      "010" when "001",
      "011" when "010",
      "000" when "011",
      "100" when "100",
      "000" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "000" when "000",
      "100" when "001",
      "000" when "010",
      "001" when "011",
      "010" when "100",
      "011" when "101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "1" when "011",
      "0" when "100",
      "0" when "101",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "1" when "011",
      "0" when "100",
      "0" when "101",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "1" when "010",
      "0" when "011",
      "0" when "100",
      "0" when "101",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1 is
signal t_in : std_logic_vector(2 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   with t_in select t_out <= 
      "0" when "000",
      "0" when "001",
      "0" when "010",
      "1" when "011",
      "0" when "100",
      "0" when "101",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(2 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
   instLUT: GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_6_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(2 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_6_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(2 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount61_out : std_logic_vector(2 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add5_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add5_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add5_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add15_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add19_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add19_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add19_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add115_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add115_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add115_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add116_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add116_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add116_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add116_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add117_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add117_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add29_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add29_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add29_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add36_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add36_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add36_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add126_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add126_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add126_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add126_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add126_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add126_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add37_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add37_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add37_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add38_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add38_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add38_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add38_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add38_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract5_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract6_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract6_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product9_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product9_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract7_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract7_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No376_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No377_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No378_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No379_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No380_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No381_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No382_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No383_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No384_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No385_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No386_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No387_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add50_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add50_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No388_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add50_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No389_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No390_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No391_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No392_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No393_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No394_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No395_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No396_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No397_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product18_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No398_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product18_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No399_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No400_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No401_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No402_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No403_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No404_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No406_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No407_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product19_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product19_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No409_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No411_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No414_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No416_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product28_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No418_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product28_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No419_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No421_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No422_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No423_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No424_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No425_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No426_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No427_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product38_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No428_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product38_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No429_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No430_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No431_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add52_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No432_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No433_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add52_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No434_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No435_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add52_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No436_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No437_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add52_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No438_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add52_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No439_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add54_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add54_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add54_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No444_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No448_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No449_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No450_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No451_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No452_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No453_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No454_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No455_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No456_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No457_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No458_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No459_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No460_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No461_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No462_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No463_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No464_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No465_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No466_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No467_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No468_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No469_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No470_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No471_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No472_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No473_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No474_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No475_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No476_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No477_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No478_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No479_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No480_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No481_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No482_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No483_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No484_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No485_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract14_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract14_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No486_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract14_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No487_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No488_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No489_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract17_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No490_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract17_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No491_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No492_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No493_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No494_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No495_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No496_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No497_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract19_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract19_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No498_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract19_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No499_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No500_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No501_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No502_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No503_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No504_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No505_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No506_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No507_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No508_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No509_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No510_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No511_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No512_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No513_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No514_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No515_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract21_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No516_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No517_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add63_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add63_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No518_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add63_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No519_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No520_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No521_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No522_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No523_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No524_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No525_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No526_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No527_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product50_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No528_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product50_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No529_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No530_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No531_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No532_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No533_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No534_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No535_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No536_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No537_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No538_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No539_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No540_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No541_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No542_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No543_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No544_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No545_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No546_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No547_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No548_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No549_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No550_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No551_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No552_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No553_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No554_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No555_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No556_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No557_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No558_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No559_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No560_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No561_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No562_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No563_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No564_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No565_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No566_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No567_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No568_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No569_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product124_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No570_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product124_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No571_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No572_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No573_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No574_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No575_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No576_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No577_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No578_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No579_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No580_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No581_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No582_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No583_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No584_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No585_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No586_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No587_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No588_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No589_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No590_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No591_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No592_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No593_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No594_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No595_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No596_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No597_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No598_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No599_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No600_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No601_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No602_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No603_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No604_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No605_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No606_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No607_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No608_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No609_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No610_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No611_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No612_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No613_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No614_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No615_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No616_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No617_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No618_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No619_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No620_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No621_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No622_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No623_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No624_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No625_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No626_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No627_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No628_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No629_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No630_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No631_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No632_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No633_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No634_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No635_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No636_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No637_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No638_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No639_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No640_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No641_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract27_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No642_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No643_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract27_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No644_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No645_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract27_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No646_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No647_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract27_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No648_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No649_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract27_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No650_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract27_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No651_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No652_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No653_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No654_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No655_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No656_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No657_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No658_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No659_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract42_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No660_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract42_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No661_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add84_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add84_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No662_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add84_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No663_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No664_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No665_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No666_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No667_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No668_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No669_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No670_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No671_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract44_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No672_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract44_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No673_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract45_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No674_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract45_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No675_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No676_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No677_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No678_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No679_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No680_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No681_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No682_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No683_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No684_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No685_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract47_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No686_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No687_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract47_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No688_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No689_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract47_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No690_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No691_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract52_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No692_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No693_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract52_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No694_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No695_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract52_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No696_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No697_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract52_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No698_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No699_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract52_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No700_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract52_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No701_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract112_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No702_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No703_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract112_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No704_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No705_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract112_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No706_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No707_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract112_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No708_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No709_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract112_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No710_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract112_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No711_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract56_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No712_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No713_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract56_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No714_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No715_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract56_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No716_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No717_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract56_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No718_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract56_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No719_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract60_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract60_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No720_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract60_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No721_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract60_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract60_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No722_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract60_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No723_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract126_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract126_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No724_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract126_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No725_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract135_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract135_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No726_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract135_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No727_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No320_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No321_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No325_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No326_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No327_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No328_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No329_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Add84_4_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add84_4_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract135_4_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract135_4_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No232_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No233_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add5_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add5_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No230_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add5_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add5_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No231_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add15_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add15_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add7_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add7_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add7_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add7_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add7_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add7_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No34_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No40_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add16_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add16_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add16_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add16_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add16_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add16_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No30_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No46_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add9_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add9_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Add9_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Add9_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No59_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No64_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No31_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Add18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Add18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No32_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Add18_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Add18_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No33_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Add19_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Add19_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Add19_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Add19_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Add115_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Add115_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Add116_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Add116_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No55_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No60_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Add116_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Add116_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No56_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No61_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Add116_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Add116_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Add117_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Add117_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Add117_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Add117_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Add117_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Add117_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No57_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No62_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Add117_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Add117_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Add29_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Add29_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No58_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No63_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Add36_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Add36_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No79_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No84_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Add126_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Add126_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No75_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No80_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Add126_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Add126_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Add37_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Add37_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No322_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No327_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Add127_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Add127_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No76_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No321_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No81_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No326_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Add127_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Add127_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No77_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No82_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Add127_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Add127_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No323_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No328_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Add38_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Add38_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No320_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No325_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Add38_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Add38_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Add38_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Add38_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Add38_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Add38_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No78_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No83_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Add128_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Add128_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Add128_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Add128_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Add128_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Add128_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No324_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No329_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Add129_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Add129_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No90_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No95_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Add129_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Add129_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No91_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No96_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Add129_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Add129_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No92_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No97_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Add129_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Add129_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Add129_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Add129_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No94_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No99_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No200_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No205_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No201_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No206_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Add40_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Add40_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No202_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No207_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Add40_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Add40_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No93_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No98_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Add40_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Add40_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Add130_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Add130_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Add130_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Add130_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Add130_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Add130_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Add130_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Add130_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No203_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No208_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Add130_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Add130_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No204_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No209_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No54_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No69_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No35_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No50_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No51_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Subtract3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Subtract3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No52_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Product13_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Product13_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Product13_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Product13_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Product13_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Product13_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Product13_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Product13_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out_to_Product13_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out_to_Product13_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No36_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No37_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No38_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No53_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out_to_Subtract6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out_to_Subtract6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No50_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No65_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out_to_Subtract6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out_to_Subtract6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No51_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No66_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out_to_Subtract6_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out_to_Subtract6_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No52_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No67_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out_to_Subtract6_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out_to_Subtract6_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No53_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No68_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out_to_Product9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out_to_Product9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out_to_Product9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out_to_Product9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out_to_Product9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out_to_Product9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out_to_Product9_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out_to_Product9_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out_to_Product9_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out_to_Product9_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out_to_Product26_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out_to_Product26_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out_to_Product26_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out_to_Product26_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out_to_Subtract7_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out_to_Subtract7_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out_to_Subtract7_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out_to_Subtract7_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out_to_Subtract7_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out_to_Subtract7_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out_to_Subtract7_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out_to_Subtract7_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out_to_Subtract7_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out_to_Subtract7_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No74_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No89_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out_to_Product17_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out_to_Product17_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out_to_Product17_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out_to_Product17_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out_to_Product17_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out_to_Product17_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out_to_Product17_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out_to_Product17_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out_to_Product17_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out_to_Product17_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No376_out_to_Product37_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No377_out_to_Product37_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No378_out_to_Product37_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No379_out_to_Product37_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No380_out_to_Product37_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No381_out_to_Product37_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No382_out_to_Product37_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No383_out_to_Product37_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No384_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No385_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No386_out_to_Subtract8_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No387_out_to_Subtract8_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No39_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No388_out_to_Add50_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No389_out_to_Add50_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No390_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No391_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No392_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No393_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No394_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No395_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No396_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No397_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No398_out_to_Product18_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No399_out_to_Product18_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No400_out_to_Product19_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No401_out_to_Product19_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No402_out_to_Product19_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No403_out_to_Product19_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No404_out_to_Product19_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No405_out_to_Product19_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No406_out_to_Product19_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No407_out_to_Product19_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No408_out_to_Product19_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No409_out_to_Product19_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No410_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No411_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No412_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No413_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No414_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No415_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No416_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No417_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No418_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No419_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No420_out_to_Product38_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No421_out_to_Product38_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No422_out_to_Product38_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No423_out_to_Product38_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No424_out_to_Product38_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No425_out_to_Product38_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No426_out_to_Product38_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No427_out_to_Product38_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No428_out_to_Product38_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No429_out_to_Product38_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No430_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No431_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No432_out_to_Add52_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No433_out_to_Add52_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No434_out_to_Add52_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No435_out_to_Add52_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No436_out_to_Add52_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No437_out_to_Add52_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No438_out_to_Add52_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No439_out_to_Add52_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No440_out_to_Add54_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No441_out_to_Add54_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No442_out_to_Add54_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No443_out_to_Add54_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No444_out_to_Add54_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No445_out_to_Add54_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No446_out_to_Product42_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No447_out_to_Product42_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No448_out_to_Product42_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No449_out_to_Product42_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No450_out_to_Product42_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No451_out_to_Product42_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No452_out_to_Product42_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No453_out_to_Product42_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No454_out_to_Product42_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No455_out_to_Product42_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No456_out_to_Product114_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No457_out_to_Product114_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No458_out_to_Product114_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No459_out_to_Product114_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No460_out_to_Product114_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No461_out_to_Product114_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No462_out_to_Product114_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No463_out_to_Product114_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No464_out_to_Product114_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No465_out_to_Product114_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No466_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No467_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No468_out_to_Product213_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No469_out_to_Product213_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No470_out_to_Product213_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No471_out_to_Product213_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No472_out_to_Product213_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No473_out_to_Product213_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No474_out_to_Product213_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No475_out_to_Product213_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No476_out_to_Product313_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No477_out_to_Product313_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No478_out_to_Product313_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No479_out_to_Product313_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No480_out_to_Product313_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No481_out_to_Product313_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No482_out_to_Product313_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No483_out_to_Product313_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No484_out_to_Product313_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No485_out_to_Product313_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No486_out_to_Subtract14_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No487_out_to_Subtract14_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No149_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No154_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No488_out_to_Subtract17_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No489_out_to_Subtract17_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No70_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No145_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No85_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No150_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No490_out_to_Subtract17_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No491_out_to_Subtract17_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No146_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No71_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No151_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No86_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No492_out_to_Subtract18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No493_out_to_Subtract18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No494_out_to_Subtract18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No495_out_to_Subtract18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No496_out_to_Subtract18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No497_out_to_Subtract18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No147_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No72_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No152_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No87_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No498_out_to_Subtract19_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No499_out_to_Subtract19_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No148_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No73_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No153_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No88_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No500_out_to_Subtract20_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No501_out_to_Subtract20_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No195_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No210_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No502_out_to_Subtract20_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No503_out_to_Subtract20_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No196_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No211_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No504_out_to_Subtract20_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No505_out_to_Subtract20_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No506_out_to_Subtract20_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No507_out_to_Subtract20_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No508_out_to_Subtract21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No509_out_to_Subtract21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No510_out_to_Subtract21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No511_out_to_Subtract21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No512_out_to_Subtract21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No513_out_to_Subtract21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No197_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No212_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No514_out_to_Subtract21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No515_out_to_Subtract21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No516_out_to_Subtract21_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No517_out_to_Subtract21_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No199_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No214_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No518_out_to_Add63_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No519_out_to_Add63_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No234_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No520_out_to_Product50_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No521_out_to_Product50_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No522_out_to_Product50_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No523_out_to_Product50_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No524_out_to_Product50_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No525_out_to_Product50_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No526_out_to_Product50_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No527_out_to_Product50_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No528_out_to_Product50_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No529_out_to_Product50_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No530_out_to_Product122_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No531_out_to_Product122_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No532_out_to_Product122_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No533_out_to_Product122_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No534_out_to_Product122_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No535_out_to_Product122_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No536_out_to_Product122_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No537_out_to_Product122_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No538_out_to_Product122_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No539_out_to_Product122_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No540_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No541_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No542_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No543_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No544_out_to_Product221_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No545_out_to_Product221_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No546_out_to_Product221_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No547_out_to_Product221_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No548_out_to_Product221_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No549_out_to_Product221_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No550_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No551_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No552_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No553_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No554_out_to_Product321_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No555_out_to_Product321_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No556_out_to_Product321_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No557_out_to_Product321_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No558_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No559_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No560_out_to_Subtract23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No561_out_to_Subtract23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No562_out_to_Product124_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No563_out_to_Product124_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No564_out_to_Product124_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No565_out_to_Product124_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No566_out_to_Product124_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No567_out_to_Product124_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No568_out_to_Product124_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No569_out_to_Product124_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No570_out_to_Product124_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No571_out_to_Product124_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No572_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No573_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No574_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No575_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No576_out_to_Product323_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No577_out_to_Product323_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No578_out_to_Product323_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No579_out_to_Product323_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No580_out_to_Product323_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No581_out_to_Product323_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No582_out_to_Subtract24_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No583_out_to_Subtract24_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No215_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No220_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No584_out_to_Subtract24_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No585_out_to_Subtract24_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No216_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No221_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No586_out_to_Subtract24_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No587_out_to_Subtract24_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No588_out_to_Subtract24_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No589_out_to_Subtract24_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No198_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No213_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No590_out_to_Subtract24_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No591_out_to_Subtract24_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No592_out_to_Subtract26_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No593_out_to_Subtract26_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No594_out_to_Subtract26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No595_out_to_Subtract26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No596_out_to_Subtract26_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No597_out_to_Subtract26_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No217_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No222_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No598_out_to_Subtract26_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No599_out_to_Subtract26_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No600_out_to_Subtract26_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No601_out_to_Subtract26_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No219_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No224_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No602_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No603_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No604_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No605_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No606_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No607_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No608_out_to_Product55_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No609_out_to_Product55_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No610_out_to_Product55_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No611_out_to_Product55_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No612_out_to_Product127_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No613_out_to_Product127_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No614_out_to_Product127_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No615_out_to_Product127_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No616_out_to_Product127_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No617_out_to_Product127_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No618_out_to_Product127_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No619_out_to_Product127_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No620_out_to_Product127_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No621_out_to_Product127_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No622_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No623_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No624_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No625_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No626_out_to_Product226_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No627_out_to_Product226_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No628_out_to_Product226_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No629_out_to_Product226_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No630_out_to_Product226_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No631_out_to_Product226_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No632_out_to_Product326_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No633_out_to_Product326_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No634_out_to_Product326_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No635_out_to_Product326_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No636_out_to_Product326_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No637_out_to_Product326_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No638_out_to_Product326_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No639_out_to_Product326_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No640_out_to_Product326_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No641_out_to_Product326_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No642_out_to_Subtract27_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No643_out_to_Subtract27_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No644_out_to_Subtract27_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No645_out_to_Subtract27_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No646_out_to_Subtract27_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No647_out_to_Subtract27_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No648_out_to_Subtract27_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No649_out_to_Subtract27_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No218_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No223_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No650_out_to_Subtract27_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No651_out_to_Subtract27_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No652_out_to_Subtract42_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No653_out_to_Subtract42_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No654_out_to_Subtract42_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No655_out_to_Subtract42_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No656_out_to_Subtract42_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No657_out_to_Subtract42_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No658_out_to_Subtract42_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No659_out_to_Subtract42_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No660_out_to_Subtract42_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No661_out_to_Subtract42_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No662_out_to_Add84_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No663_out_to_Add84_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Add84_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Add84_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Add84_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Add84_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No664_out_to_Subtract44_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No665_out_to_Subtract44_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No666_out_to_Subtract44_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No667_out_to_Subtract44_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No668_out_to_Subtract44_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No669_out_to_Subtract44_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No670_out_to_Subtract44_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No671_out_to_Subtract44_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No672_out_to_Subtract44_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No673_out_to_Subtract44_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No674_out_to_Subtract45_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No675_out_to_Subtract45_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No676_out_to_Subtract46_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No677_out_to_Subtract46_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No235_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No678_out_to_Subtract46_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No679_out_to_Subtract46_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No236_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No680_out_to_Subtract46_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No681_out_to_Subtract46_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No237_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No682_out_to_Subtract46_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No683_out_to_Subtract46_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No238_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No684_out_to_Subtract46_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No685_out_to_Subtract46_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No239_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No686_out_to_Subtract47_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No687_out_to_Subtract47_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No688_out_to_Subtract47_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No689_out_to_Subtract47_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No690_out_to_Subtract47_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No691_out_to_Subtract47_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No134_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No692_out_to_Subtract52_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No693_out_to_Subtract52_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No694_out_to_Subtract52_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No695_out_to_Subtract52_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No696_out_to_Subtract52_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No697_out_to_Subtract52_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No698_out_to_Subtract52_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No699_out_to_Subtract52_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No700_out_to_Subtract52_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No701_out_to_Subtract52_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No702_out_to_Subtract112_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No703_out_to_Subtract112_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No704_out_to_Subtract112_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No705_out_to_Subtract112_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No706_out_to_Subtract112_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No707_out_to_Subtract112_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No708_out_to_Subtract112_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No709_out_to_Subtract112_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No710_out_to_Subtract112_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No711_out_to_Subtract112_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No712_out_to_Subtract56_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No713_out_to_Subtract56_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No714_out_to_Subtract56_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No715_out_to_Subtract56_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No716_out_to_Subtract56_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No717_out_to_Subtract56_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No718_out_to_Subtract56_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No719_out_to_Subtract56_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No720_out_to_Subtract60_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No721_out_to_Subtract60_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No722_out_to_Subtract60_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No723_out_to_Subtract60_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No724_out_to_Subtract126_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No725_out_to_Subtract126_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No54_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No726_out_to_Subtract135_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No727_out_to_Subtract135_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract135_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Subtract135_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Subtract135_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract135_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount61_instance: ModuloCounter_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount61_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg119_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg119_out;
SharedReg136_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg136_out;
SharedReg139_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg142_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg142_out;
SharedReg116_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg119_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg136_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg139_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg142_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg133_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg158_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg158_out;
SharedReg167_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg167_out;
SharedReg179_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg179_out;
SharedReg130_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg130_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg158_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg167_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg179_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg130_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg75_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg66_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg55_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg70_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg70_out;
SharedReg94_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg94_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg70_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg94_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg99_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg77_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg68_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg81_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg81_out;
SharedReg96_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg96_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg81_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg96_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg63_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg66_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg68_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg81_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg81_out;
SharedReg72_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg72_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg81_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg72_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg75_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg77_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg79_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg101_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg83_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg83_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg79_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg83_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg133_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg136_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg136_out;
SharedReg125_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg127_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg130_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg130_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg136_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg125_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg127_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg130_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg161_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg158_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg158_out;
SharedReg139_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg142_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg142_out;
SharedReg145_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg145_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg158_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg139_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg142_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg145_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg161_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg161_out;
SharedReg164_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg164_out;
SharedReg177_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg177_out;
SharedReg182_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg182_out;
SharedReg145_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg145_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg161_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg164_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg177_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg182_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg145_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg49_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg52_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg52_out;
SharedReg55_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg70_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg70_out;
SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg60_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg52_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg70_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg60_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg106_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg109_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg109_out;
SharedReg79_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg101_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg103_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg103_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg109_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg79_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg103_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg119_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg119_out;
SharedReg122_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg122_out;
SharedReg111_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg111_out;
SharedReg114_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg116_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg116_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg119_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg111_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg116_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg99_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg109_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg109_out;
SharedReg111_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg111_out;
SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg94_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg94_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg109_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg111_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg94_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg106_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg122_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg122_out;
SharedReg125_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg127_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg127_out;
SharedReg96_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg96_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg125_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg127_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg96_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg171_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg171_out;
SharedReg164_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg164_out;
SharedReg167_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg167_out;
SharedReg179_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg179_out;
SharedReg185_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg185_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg171_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg164_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg167_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg179_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg185_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg188_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg188_out;
SharedReg174_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg174_out;
SharedReg177_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg177_out;
SharedReg182_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg182_out;
SharedReg191_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg191_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg188_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg177_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg182_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg191_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg849_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg851_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg851_out;
SharedReg853_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg853_out;
SharedReg855_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg895_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg895_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg851_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg853_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg895_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg893_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg893_out;
SharedReg693_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg693_out;
SharedReg520_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg520_out;
SharedReg473_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg473_out;
SharedReg897_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg897_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg893_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg693_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg520_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg473_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg897_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg865_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg865_out;
SharedReg801_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg801_out;
SharedReg803_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg803_out;
SharedReg847_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg847_out;
SharedReg873_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg873_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg865_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg801_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg803_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg847_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg873_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg875_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg875_out;
SharedReg867_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg867_out;
SharedReg858_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg858_out;
SharedReg860_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg860_out;
SharedReg883_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg883_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg875_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg867_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg858_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg860_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg883_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg798_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg798_out;
SharedReg801_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg801_out;
SharedReg858_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg858_out;
SharedReg860_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg860_out;
SharedReg808_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg808_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg798_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg801_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg858_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg860_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg808_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg865_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg865_out;
SharedReg867_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg867_out;
SharedReg869_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg869_out;
SharedReg871_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg871_out;
SharedReg862_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg862_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg865_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg867_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg869_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg871_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg862_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg828_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg828_out;
SharedReg814_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg814_out;
SharedReg889_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg889_out;
SharedReg891_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg891_out;
SharedReg856_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg856_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg828_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg814_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg889_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg891_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg856_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg849_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg832_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg832_out;
SharedReg817_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg817_out;
SharedReg820_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg820_out;
SharedReg895_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg895_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg832_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg817_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg820_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg895_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg354_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg354_out;
SharedReg357_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg360_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg360_out;
SharedReg397_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg397_out;
SharedReg897_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg897_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg354_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg360_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg897_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg738_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg738_out;
SharedReg742_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg742_out;
SharedReg803_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg803_out;
SharedReg847_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg847_out;
SharedReg754_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg754_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg738_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg742_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg803_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg847_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg754_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg885_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg885_out;
SharedReg877_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg877_out;
SharedReg869_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg869_out;
SharedReg871_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg871_out;
SharedReg824_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg824_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg885_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg877_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg869_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg871_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg824_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg811_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg811_out;
SharedReg887_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg887_out;
SharedReg879_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg879_out;
SharedReg881_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg881_out;
SharedReg843_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg843_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg811_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg887_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg879_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg881_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg843_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg875_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg875_out;
SharedReg877_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg877_out;
SharedReg879_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg879_out;
SharedReg881_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg881_out;
SharedReg873_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg873_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg875_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg877_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg879_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg881_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg873_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg885_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg885_out;
SharedReg887_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg887_out;
SharedReg889_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg889_out;
SharedReg891_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg891_out;
SharedReg883_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg883_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg885_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg887_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg889_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg891_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg883_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg893_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg893_out;
SharedReg851_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg851_out;
SharedReg836_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg836_out;
SharedReg840_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg840_out;
SharedReg897_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg897_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg893_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg851_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg836_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg840_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg897_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg354_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg354_out;
SharedReg693_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg693_out;
SharedReg853_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg853_out;
SharedReg855_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg898_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg898_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg354_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg693_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg853_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg898_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg638_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg638_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg607_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg607_out;
SharedReg190_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg190_out;
SharedReg606_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg606_out;
SharedReg246_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg246_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg638_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg607_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg190_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg606_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg246_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg353_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg799_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg799_out;
SharedReg224_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg798_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg798_out;
SharedReg119_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg119_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg799_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg798_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg119_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg228_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg228_out;
SharedReg643_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg643_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg_out;
SharedReg611_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg611_out;
SharedReg200_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg200_out;
SharedReg247_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg247_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg228_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg643_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg611_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg200_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg247_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg136_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg356_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg356_out;
SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg802_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg802_out;
SharedReg215_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg215_out;
SharedReg148_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg148_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg356_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg802_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg215_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg148_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg250_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg250_out;
SharedReg233_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg233_out;
SharedReg649_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg649_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg_out;
SharedReg389_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg389_out;
SharedReg443_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg443_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg250_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg233_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg649_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg389_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg443_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg153_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg139_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg695_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg695_out;
SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg16_out;
SharedReg629_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg629_out;
SharedReg747_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg747_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg695_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg629_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg747_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg206_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg650_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg650_out;
Delay3No232_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= Delay3No232_out;
SharedReg677_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg677_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg362_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg362_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg650_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No232_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg677_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg362_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg207_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg860_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg860_out;
SharedReg792_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg792_out;
SharedReg685_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg685_out;
SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg618_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg618_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg860_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg792_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg685_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg618_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg596_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg596_out;
SharedReg774_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg774_out;
SharedReg670_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg670_out;
SharedReg679_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg679_out;
SharedReg658_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg658_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg596_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg774_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg670_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg679_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg658_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg809_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg809_out;
SharedReg784_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg784_out;
SharedReg774_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg774_out;
SharedReg686_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg686_out;
SharedReg400_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg400_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg809_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg784_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg774_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg686_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg245_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg245_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg352_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg352_out;
SharedReg210_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg210_out;
SharedReg244_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg244_out;
SharedReg436_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg436_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg245_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg352_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg210_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg244_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg436_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No42_out);

SharedReg261_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg621_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg621_out;
SharedReg211_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg211_out;
SharedReg538_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg538_out;
SharedReg849_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg849_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg621_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg211_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg538_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg849_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg407_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg407_out;
SharedReg248_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg248_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg385_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg385_out;
SharedReg604_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg604_out;
SharedReg439_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg439_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg407_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg248_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg385_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg604_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg439_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No44_out);

SharedReg851_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg851_out;
SharedReg264_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
SharedReg625_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg625_out;
SharedReg744_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg744_out;
SharedReg405_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg405_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg851_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg625_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg744_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg405_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg442_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg442_out;
SharedReg410_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg410_out;
SharedReg251_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg251_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1_out;
SharedReg532_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg532_out;
SharedReg358_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg358_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg442_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg410_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg251_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg532_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg358_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No46_out);

SharedReg408_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg408_out;
SharedReg853_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg853_out;
SharedReg267_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg267_out;
SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg265_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg648_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg648_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg408_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg853_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg267_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg648_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg413_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg413_out;
SharedReg268_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg268_out;
SharedReg254_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg254_out;
SharedReg653_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg653_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg536_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg536_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg413_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg268_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg254_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg653_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg536_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No48_out);

SharedReg751_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg751_out;
SharedReg45_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg45_out;
SharedReg142_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg521_out;
SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg17_out;
SharedReg269_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg269_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg751_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg45_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg521_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg269_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg474_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg474_out;
SharedReg187_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg187_out;
Delay3No233_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= Delay3No233_out;
SharedReg288_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg288_out;
SharedReg258_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg258_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg474_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg187_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No233_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg288_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg258_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No50_out);

SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg17_out;
SharedReg633_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg633_out;
SharedReg258_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg258_out;
SharedReg794_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg103_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg103_out;
SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg273_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg633_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg258_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg794_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg103_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_0_impl_out,
                 X => Delay1No52_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg403_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg403_out;
SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg524_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg524_out;
SharedReg601_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg601_out;
SharedReg600_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg600_out;
SharedReg276_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg276_out;
   MUX_Add3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg403_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg524_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg601_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg600_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg276_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_0_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_0_out,
                 Y => Delay1No52_out);

SharedReg437_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg437_out;
SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg275_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg275_out;
SharedReg740_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg740_out;
SharedReg402_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg402_out;
SharedReg86_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg86_out;
   MUX_Add3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg437_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg275_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg740_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg402_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg86_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_0_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_1_impl_out,
                 X => Delay1No54_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg263_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg263_out;
SharedReg406_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg406_out;
SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg528_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg528_out;
SharedReg384_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg384_out;
SharedReg279_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg279_out;
   MUX_Add3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg263_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg406_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg528_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg384_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg279_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_1_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_0_out,
                 Y => Delay1No54_out);

SharedReg90_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg440_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg440_out;
SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg18_out;
SharedReg279_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg279_out;
SharedReg627_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg213_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg213_out;
   MUX_Add3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg440_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg279_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg213_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_1_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_2_impl_out,
                 X => Delay1No56_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast);

SharedReg282_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg282_out;
SharedReg266_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg266_out;
SharedReg409_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg409_out;
SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg2_out;
SharedReg410_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg410_out;
SharedReg251_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg251_out;
   MUX_Add3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg266_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg409_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg410_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg251_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_2_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_0_out,
                 Y => Delay1No56_out);

SharedReg217_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg217_out;
SharedReg41_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg445_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg445_out;
SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg18_out;
SharedReg727_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg727_out;
SharedReg235_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg235_out;
   MUX_Add3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg217_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg445_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg727_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg235_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_2_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add3_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_3_impl_out,
                 X => Delay1No58_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg361_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg361_out;
SharedReg447_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg447_out;
SharedReg413_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg269_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg269_out;
SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg330_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg330_out;
   MUX_Add3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg361_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg447_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg413_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg269_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg330_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_3_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_0_out,
                 Y => Delay1No58_out);

SharedReg733_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg733_out;
SharedReg411_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg411_out;
SharedReg855_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg855_out;
SharedReg286_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg286_out;
SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg731_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg731_out;
   MUX_Add3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg733_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg411_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg855_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg286_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg731_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_3_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add3_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_4_impl_out,
                 X => Delay1No60_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast);

SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg2_out;
SharedReg478_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg478_out;
SharedReg242_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg242_out;
SharedReg632_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg632_out;
SharedReg597_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg597_out;
SharedReg333_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg333_out;
   MUX_Add3_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg478_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg242_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg632_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg597_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg333_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_4_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_0_out,
                 Y => Delay1No60_out);

SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg287_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg287_out;
SharedReg193_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg193_out;
SharedReg862_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg862_out;
SharedReg856_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg856_out;
SharedReg396_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg396_out;
   MUX_Add3_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg287_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg193_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg862_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg856_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add3_4_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_0_impl_out,
                 X => Delay1No62_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg162_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg162_out;
SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg404_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg317_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg317_out;
SharedReg523_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg523_out;
SharedReg318_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg318_out;
   MUX_Add12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg162_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg317_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg523_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg318_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_0_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_0_out,
                 Y => Delay1No62_out);

SharedReg173_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg173_out;
SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg717_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg717_out;
SharedReg623_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg623_out;
SharedReg209_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg209_out;
SharedReg350_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg350_out;
   MUX_Add12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg173_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg717_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg623_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg209_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_0_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_1_impl_out,
                 X => Delay1No64_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg385_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg385_out;
SharedReg165_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg407_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg262_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg262_out;
SharedReg603_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg603_out;
   MUX_Add12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg385_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg262_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg603_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_1_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_0_out,
                 Y => Delay1No64_out);

SharedReg383_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg383_out;
SharedReg176_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg176_out;
SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg722_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg230_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg230_out;
SharedReg438_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg438_out;
   MUX_Add12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg383_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg230_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg438_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_1_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_2_impl_out,
                 X => Delay1No66_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg615_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg615_out;
SharedReg389_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg178_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg178_out;
SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg43_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg43_out;
SharedReg388_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg388_out;
   MUX_Add12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg615_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg178_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg43_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg388_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_2_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_0_out,
                 Y => Delay1No66_out);

SharedReg441_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg441_out;
SharedReg387_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg387_out;
SharedReg198_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg19_out;
SharedReg282_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg282_out;
SharedReg748_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg748_out;
   MUX_Add12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg441_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg387_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg198_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg282_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg748_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_2_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_3_impl_out,
                 X => Delay1No68_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg269_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg269_out;
SharedReg535_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg535_out;
SharedReg285_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg285_out;
SharedReg412_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg412_out;
SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg47_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg47_out;
   MUX_Add12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg269_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg535_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg285_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg412_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg47_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_3_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_0_out,
                 Y => Delay1No68_out);

SharedReg256_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg236_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg236_out;
SharedReg60_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg60_out;
SharedReg449_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg449_out;
SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg19_out;
SharedReg284_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg284_out;
   MUX_Add12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg236_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg60_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg449_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg284_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_3_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_4_impl_out,
                 X => Delay1No70_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg334_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg334_out;
SharedReg452_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg452_out;
SharedReg270_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg270_out;
SharedReg548_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg131_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg131_out;
   MUX_Add12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg334_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg452_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg270_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg131_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_4_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_0_out,
                 Y => Delay1No70_out);

SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg735_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg735_out;
SharedReg756_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg660_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg660_out;
SharedReg660_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg660_out;
SharedReg147_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
   MUX_Add12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg735_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg756_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg660_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg660_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg147_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add12_4_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add5_1_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add5_1_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add5_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add5_1_impl_out,
                 X => Delay1No72_out_to_Add5_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add5_1_impl_parent_implementedSystem_port_1_cast);

Delay3No230_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No230_out;
SharedReg673_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg673_out;
SharedReg769_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg769_out;
SharedReg779_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg779_out;
SharedReg201_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg201_out;
SharedReg610_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg610_out;
   MUX_Add5_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No230_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg673_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg769_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg779_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg201_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg610_out_to_MUX_Add5_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add5_1_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_1_impl_0_out,
                 Y => Delay1No72_out);

SharedReg788_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg788_out;
SharedReg683_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg683_out;
SharedReg779_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg779_out;
SharedReg788_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg788_out;
SharedReg214_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg214_out;
SharedReg801_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg801_out;
   MUX_Add5_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg788_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg683_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg779_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg788_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg214_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg801_out_to_MUX_Add5_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add5_1_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_1_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add5_2_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add5_2_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add5_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add5_2_impl_out,
                 X => Delay1No74_out_to_Add5_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add5_2_impl_parent_implementedSystem_port_1_cast);

SharedReg628_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg628_out;
Delay3No231_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_2_cast <= Delay3No231_out;
SharedReg675_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg675_out;
SharedReg771_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg771_out;
SharedReg615_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg615_out;
SharedReg196_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg196_out;
   MUX_Add5_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg628_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No231_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg675_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg771_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg615_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg196_out_to_MUX_Add5_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add5_2_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_2_impl_0_out,
                 Y => Delay1No74_out);

SharedReg858_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg858_out;
SharedReg790_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg790_out;
SharedReg684_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg684_out;
SharedReg781_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg781_out;
SharedReg804_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg804_out;
SharedReg204_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg204_out;
   MUX_Add5_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg858_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg790_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg684_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg781_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg804_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg204_out_to_MUX_Add5_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add5_2_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add5_2_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add6_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add6_4_impl_out,
                 X => Delay1No76_out_to_Add6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg4_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg662_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg662_out;
SharedReg333_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg333_out;
SharedReg633_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg633_out;
SharedReg395_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg395_out;
SharedReg451_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg451_out;
   MUX_Add6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg662_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg333_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg633_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg395_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg451_out_to_MUX_Add6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add6_4_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_4_impl_0_out,
                 Y => Delay1No76_out);

SharedReg20_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg477_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg477_out;
SharedReg635_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg635_out;
SharedReg393_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg393_out;
SharedReg473_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg473_out;
SharedReg598_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg598_out;
   MUX_Add6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg477_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg635_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg393_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg473_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg598_out_to_MUX_Add6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add6_4_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_4_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add15_4_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add15_4_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add15_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add15_4_impl_out,
                 X => Delay1No78_out_to_Add15_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add15_4_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg398_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg398_out;
SharedReg477_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg477_out;
SharedReg661_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg661_out;
SharedReg475_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg475_out;
SharedReg186_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg186_out;
   MUX_Add15_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg398_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg477_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg661_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg475_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg186_out_to_MUX_Add15_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add15_4_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_4_impl_0_out,
                 Y => Delay1No78_out);

SharedReg21_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg333_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg333_out;
SharedReg243_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg243_out;
SharedReg241_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg596_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg596_out;
SharedReg194_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg194_out;
   MUX_Add15_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg243_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg596_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg194_out_to_MUX_Add15_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add15_4_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_4_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add7_0_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add7_0_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add7_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_0_impl_out,
                 X => Delay1No80_out_to_Add7_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add7_0_impl_parent_implementedSystem_port_1_cast);

SharedReg600_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg600_out;
SharedReg4_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg88_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg275_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg275_out;
SharedReg607_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg607_out;
SharedReg353_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg353_out;
   MUX_Add7_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg600_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg275_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg607_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg353_out_to_MUX_Add7_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add7_0_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_0_impl_0_out,
                 Y => Delay1No80_out);

SharedReg609_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg20_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg523_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg523_out;
SharedReg225_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg225_out;
SharedReg434_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg434_out;
SharedReg600_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg600_out;
   MUX_Add7_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg523_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg225_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg434_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg600_out_to_MUX_Add7_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add7_0_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_0_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add7_3_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add7_3_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add7_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_3_impl_out,
                 X => Delay1No82_out_to_Add7_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add7_3_impl_parent_implementedSystem_port_1_cast);

SharedReg391_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg618_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg618_out;
SharedReg392_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg183_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg183_out;
SharedReg4_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg361_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg361_out;
   MUX_Add7_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg618_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg183_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg4_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg361_out_to_MUX_Add7_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add7_3_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_3_impl_0_out,
                 Y => Delay1No82_out);

SharedReg807_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg807_out;
SharedReg446_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg446_out;
SharedReg390_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg208_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg208_out;
SharedReg20_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg391_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg391_out;
   MUX_Add7_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg807_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg446_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg208_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg391_out_to_MUX_Add7_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add7_3_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_3_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add7_4_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add7_4_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add7_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_4_impl_out,
                 X => Delay1No84_out_to_Add7_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add7_4_impl_parent_implementedSystem_port_1_cast);

SharedReg12_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg399_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg394_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg394_out;
SharedReg656_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg656_out;
SharedReg272_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg272_out;
Delay3No34_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_6_cast <= Delay3No34_out;
   MUX_Add7_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg394_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg656_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No34_out_to_MUX_Add7_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add7_4_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_4_impl_0_out,
                 Y => Delay1No84_out);

SharedReg28_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg28_out;
SharedReg394_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg394_out;
SharedReg737_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg737_out;
SharedReg450_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg450_out;
SharedReg289_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg289_out;
SharedReg299_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg299_out;
   MUX_Add7_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg28_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg394_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg737_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg450_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg289_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg299_out_to_MUX_Add7_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add7_4_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_4_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add16_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_0_impl_out,
                 X => Delay1No86_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast);

SharedReg189_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg5_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg317_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg403_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg403_out;
SharedReg539_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg539_out;
Delay4No40_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_6_cast <= Delay4No40_out;
   MUX_Add16_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg317_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg403_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg539_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No40_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_0_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_0_impl_0_out,
                 Y => Delay1No86_out);

SharedReg212_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg212_out;
SharedReg21_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg403_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg403_out;
SharedReg720_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg720_out;
SharedReg223_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg223_out;
SharedReg260_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg260_out;
   MUX_Add16_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg212_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg403_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg720_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg223_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg260_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_0_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_0_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add16_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_1_impl_out,
                 X => Delay1No88_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast);

SharedReg386_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg386_out;
SharedReg603_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg603_out;
SharedReg4_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg4_out;
SharedReg92_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg92_out;
SharedReg321_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg321_out;
SharedReg527_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg527_out;
   MUX_Add16_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg386_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg603_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg4_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg321_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_1_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_1_impl_0_out,
                 Y => Delay1No88_out);

SharedReg603_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg603_out;
SharedReg613_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg613_out;
SharedReg20_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg527_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg527_out;
SharedReg725_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg725_out;
SharedReg226_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg226_out;
   MUX_Add16_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg603_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg613_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg527_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg725_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg226_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_1_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_1_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add16_2_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add16_2_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add16_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_2_impl_out,
                 X => Delay1No90_out_to_Add16_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add16_2_impl_parent_implementedSystem_port_1_cast);

SharedReg531_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg531_out;
SharedReg359_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg359_out;
SharedReg615_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg615_out;
SharedReg4_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg4_out;
SharedReg388_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg388_out;
SharedReg265_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg265_out;
   MUX_Add16_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg531_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg359_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg615_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg388_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg265_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_2_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_2_impl_0_out,
                 Y => Delay1No90_out);

SharedReg231_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg231_out;
SharedReg615_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg615_out;
SharedReg631_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg631_out;
SharedReg20_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg20_out;
SharedReg325_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg325_out;
SharedReg283_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg283_out;
   MUX_Add16_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg231_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg615_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg631_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg20_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg325_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg283_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_2_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_2_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add16_3_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add16_3_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add16_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_3_impl_out,
                 X => Delay1No92_out_to_Add16_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add16_3_impl_parent_implementedSystem_port_1_cast);

SharedReg284_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg284_out;
SharedReg543_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg543_out;
SharedReg521_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg521_out;
SharedReg618_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg618_out;
SharedReg5_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg392_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg392_out;
   MUX_Add16_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg284_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg543_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg521_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg618_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg392_out_to_MUX_Add16_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_3_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_3_impl_0_out,
                 Y => Delay1No92_out);

SharedReg537_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg537_out;
SharedReg252_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg252_out;
SharedReg618_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg618_out;
SharedReg654_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg654_out;
SharedReg21_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg329_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg329_out;
   MUX_Add16_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg537_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg618_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg654_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg329_out_to_MUX_Add16_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_3_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_3_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add16_4_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add16_4_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add16_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_4_impl_out,
                 X => Delay1No94_out_to_Add16_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add16_4_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg548_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg548_out;
SharedReg547_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg547_out;
SharedReg827_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg827_out;
SharedReg656_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg656_out;
SharedReg339_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg339_out;
   MUX_Add16_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg548_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg547_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg827_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg656_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg339_out_to_MUX_Add16_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_4_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_4_impl_0_out,
                 Y => Delay1No94_out);

SharedReg22_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg242_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg242_out;
SharedReg290_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg257_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg257_out;
SharedReg401_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg401_out;
SharedReg344_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg344_out;
   MUX_Add16_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg242_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg290_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg257_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg401_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg344_out_to_MUX_Add16_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add16_4_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_4_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_0_impl_out,
                 X => Delay1No96_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast);

Delay3No30_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No30_out;
SharedReg12_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg318_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg523_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg523_out;
SharedReg350_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg350_out;
SharedReg621_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg621_out;
   MUX_Add9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No30_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg318_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg523_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg350_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg621_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_0_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_0_impl_0_out,
                 Y => Delay1No96_out);

SharedReg291_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg291_out;
SharedReg28_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg435_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg435_out;
SharedReg277_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg277_out;
SharedReg403_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg403_out;
SharedReg319_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg319_out;
   MUX_Add9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg435_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg277_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg403_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg319_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_0_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_0_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_1_impl_out,
                 X => Delay1No98_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg229_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg229_out;
SharedReg200_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg200_out;
SharedReg5_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg321_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg321_out;
SharedReg279_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg279_out;
SharedReg383_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg383_out;
   MUX_Add9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg229_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg200_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg321_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg279_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg383_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_1_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_1_impl_0_out,
                 Y => Delay1No98_out);

Delay4No46_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast <= Delay4No46_out;
SharedReg216_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg216_out;
SharedReg21_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg406_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg406_out;
SharedReg280_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg280_out;
SharedReg321_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg321_out;
   MUX_Add9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No46_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg216_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg21_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg406_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg280_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg321_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_1_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_1_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add9_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_2_impl_out,
                 X => Delay1No100_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg387_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg387_out;
SharedReg219_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg219_out;
SharedReg203_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg203_out;
SharedReg5_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg326_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg325_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg325_out;
   MUX_Add9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg387_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg219_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg203_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg5_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg326_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg325_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_2_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_2_impl_0_out,
                 Y => Delay1No100_out);

SharedReg325_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg325_out;
SharedReg234_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg234_out;
SharedReg220_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg21_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
SharedReg409_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg409_out;
SharedReg819_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg819_out;
   MUX_Add9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg325_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg234_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg220_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg409_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg819_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_2_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_2_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add9_3_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add9_3_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add9_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_3_impl_out,
                 X => Delay1No102_out_to_Add9_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add9_3_impl_parent_implementedSystem_port_1_cast);

SharedReg329_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg329_out;
SharedReg390_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg390_out;
SharedReg239_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg239_out;
SharedReg222_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg222_out;
SharedReg12_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg544_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg544_out;
   MUX_Add9_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg329_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg390_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg239_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg222_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg544_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_3_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_3_impl_0_out,
                 Y => Delay1No102_out);

SharedReg823_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg823_out;
SharedReg329_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg329_out;
SharedReg255_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg255_out;
SharedReg240_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg240_out;
SharedReg28_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg222_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg222_out;
   MUX_Add9_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg823_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg329_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg255_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg240_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg222_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_3_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_3_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Add9_4_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Add9_4_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Add9_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_4_impl_out,
                 X => Delay1No104_out_to_Add9_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Add9_4_impl_parent_implementedSystem_port_1_cast);

SharedReg7_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg7_out;
SharedReg258_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg258_out;
SharedReg451_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg397_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg397_out;
SharedReg287_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg287_out;
Delay4No59_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_6_cast <= Delay4No59_out;
   MUX_Add9_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg7_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg258_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg451_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg287_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No59_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_4_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_4_impl_0_out,
                 Y => Delay1No104_out);

SharedReg23_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg547_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg547_out;
SharedReg826_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg826_out;
SharedReg451_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg451_out;
SharedReg118_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg118_out;
Delay4No64_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No64_out;
   MUX_Add9_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg547_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg826_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg451_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg118_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No64_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add9_4_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_4_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Add18_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_0_impl_out,
                 X => Delay1No106_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg335_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg335_out;
SharedReg6_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg540_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg540_out;
SharedReg435_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg435_out;
SharedReg188_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg188_out;
SharedReg259_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg259_out;
   MUX_Add18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg335_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg540_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg435_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg188_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg259_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_0_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_0_impl_0_out,
                 Y => Delay1No106_out);

SharedReg340_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg22_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg224_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg224_out;
SharedReg813_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg813_out;
SharedReg259_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg259_out;
SharedReg135_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg135_out;
   MUX_Add18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg224_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg813_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg135_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_0_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_0_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Add18_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_1_impl_out,
                 X => Delay1No108_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg625_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg625_out;
Delay3No31_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast <= Delay3No31_out;
SharedReg12_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg322_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg322_out;
SharedReg406_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg199_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg199_out;
   MUX_Add18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg625_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No31_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg12_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg322_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg199_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_1_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_1_impl_0_out,
                 Y => Delay1No108_out);

SharedReg323_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg323_out;
SharedReg293_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg293_out;
SharedReg28_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg439_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg439_out;
SharedReg816_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg816_out;
SharedReg248_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg248_out;
   MUX_Add18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg323_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg293_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg28_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg439_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg816_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg248_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_1_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_1_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Add18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Add18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Add18_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_2_impl_out,
                 X => Delay1No110_out_to_Add18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Add18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg202_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg646_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg646_out;
Delay3No32_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_3_cast <= Delay3No32_out;
SharedReg12_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg12_out;
SharedReg155_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg155_out;
SharedReg282_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg282_out;
   MUX_Add18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg646_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No32_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg12_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg155_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg282_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_2_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_2_impl_0_out,
                 Y => Delay1No110_out);

SharedReg251_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg251_out;
SharedReg327_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg327_out;
SharedReg295_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg295_out;
SharedReg28_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg28_out;
SharedReg218_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg533_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg533_out;
   MUX_Add18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg251_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg295_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg28_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg533_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_2_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_2_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Add18_3_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Add18_3_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Add18_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_3_impl_out,
                 X => Delay1No112_out_to_Add18_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Add18_3_impl_parent_implementedSystem_port_1_cast);

SharedReg535_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg535_out;
SharedReg221_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg221_out;
SharedReg731_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg731_out;
Delay3No33_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_4_cast <= Delay3No33_out;
SharedReg6_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg6_out;
SharedReg237_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg237_out;
   MUX_Add18_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg535_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg731_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No33_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg6_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg237_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_3_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_3_impl_0_out,
                 Y => Delay1No112_out);

SharedReg545_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg545_out;
SharedReg269_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg269_out;
SharedReg331_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg331_out;
SharedReg297_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg297_out;
SharedReg22_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg535_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg535_out;
   MUX_Add18_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg545_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg269_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg331_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg297_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg22_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg535_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_3_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_3_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Add18_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_4_impl_out,
                 X => Delay1No114_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast);

SharedReg8_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg271_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg271_out;
SharedReg661_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg661_out;
SharedReg191_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg755_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg755_out;
SharedReg372_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg372_out;
   MUX_Add18_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg271_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg661_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg191_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg755_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg372_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_4_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_4_impl_0_out,
                 Y => Delay1No114_out);

SharedReg24_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg661_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg661_out;
SharedReg479_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg479_out;
SharedReg477_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg477_out;
SharedReg659_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg659_out;
SharedReg377_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg377_out;
   MUX_Add18_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg661_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg479_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg477_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg659_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg377_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add18_4_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_4_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Add19_2_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Add19_2_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Add19_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add19_2_impl_out,
                 X => Delay1No116_out_to_Add19_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Add19_2_impl_parent_implementedSystem_port_1_cast);

SharedReg770_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg770_out;
SharedReg666_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg666_out;
SharedReg369_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg369_out;
SharedReg675_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg675_out;
SharedReg781_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg781_out;
SharedReg197_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg197_out;
   MUX_Add19_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg770_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg666_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg369_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg675_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg781_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Add19_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add19_2_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_2_impl_0_out,
                 Y => Delay1No116_out);

SharedReg780_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg780_out;
SharedReg770_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg770_out;
SharedReg374_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg374_out;
SharedReg684_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg684_out;
SharedReg790_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg790_out;
SharedReg203_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg203_out;
   MUX_Add19_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg780_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg770_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg374_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg684_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg790_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg203_out_to_MUX_Add19_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add19_2_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_2_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Add19_3_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Add19_3_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Add19_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add19_3_impl_out,
                 X => Delay1No118_out_to_Add19_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Add19_3_impl_parent_implementedSystem_port_1_cast);

SharedReg184_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg772_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg772_out;
SharedReg668_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg668_out;
SharedReg370_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg370_out;
SharedReg773_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg773_out;
SharedReg447_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg447_out;
   MUX_Add19_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg772_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg668_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg370_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg773_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg447_out_to_MUX_Add19_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add19_3_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_3_impl_0_out,
                 Y => Delay1No118_out);

SharedReg222_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg222_out;
SharedReg782_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg782_out;
SharedReg772_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg772_out;
SharedReg375_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg375_out;
SharedReg783_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg783_out;
SharedReg805_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg805_out;
   MUX_Add19_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg222_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg782_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg772_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg375_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg783_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg805_out_to_MUX_Add19_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add19_3_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add19_3_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Add115_1_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Add115_1_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Add115_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add115_1_impl_out,
                 X => Delay1No120_out_to_Add115_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Add115_1_impl_parent_implementedSystem_port_1_cast);

SharedReg262_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg336_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg336_out;
SharedReg6_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg150_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg150_out;
SharedReg527_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg527_out;
SharedReg320_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg320_out;
   MUX_Add115_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg6_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg150_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg527_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg320_out_to_MUX_Add115_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add115_1_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add115_1_impl_0_out,
                 Y => Delay1No120_out);

SharedReg160_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg341_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg341_out;
SharedReg22_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg227_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg227_out;
SharedReg529_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg529_out;
SharedReg640_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg640_out;
   MUX_Add115_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg22_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg227_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg529_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg640_out_to_MUX_Add115_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add115_1_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add115_1_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Add116_0_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Add116_0_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Add116_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add116_0_impl_out,
                 X => Delay1No122_out_to_Add116_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Add116_0_impl_parent_implementedSystem_port_1_cast);

Delay4No55_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No55_out;
SharedReg7_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg245_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg539_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg539_out;
SharedReg316_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg316_out;
SharedReg717_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg717_out;
   MUX_Add116_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No55_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg245_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg539_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg316_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg717_out_to_MUX_Add116_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add116_0_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_0_impl_0_out,
                 Y => Delay1No122_out);

Delay4No60_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No60_out;
SharedReg23_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg539_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg539_out;
SharedReg525_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg525_out;
SharedReg636_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg636_out;
SharedReg639_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg639_out;
   MUX_Add116_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No60_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg539_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg525_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg636_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg639_out_to_MUX_Add116_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add116_0_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_0_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Add116_1_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Add116_1_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Add116_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add116_1_impl_out,
                 X => Delay1No124_out_to_Add116_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Add116_1_impl_parent_implementedSystem_port_1_cast);

SharedReg722_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg722_out;
Delay4No56_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No56_out;
SharedReg7_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg7_out;
SharedReg248_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg248_out;
SharedReg439_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg439_out;
SharedReg174_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg174_out;
   MUX_Add116_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg722_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No56_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg7_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg248_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg439_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg174_out_to_MUX_Add116_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add116_1_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_1_impl_0_out,
                 Y => Delay1No124_out);

SharedReg644_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg644_out;
Delay4No61_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No61_out;
SharedReg23_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg149_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg149_out;
SharedReg835_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg278_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg278_out;
   MUX_Add116_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg644_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No61_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg23_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg149_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg278_out_to_MUX_Add116_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add116_1_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_1_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Add116_2_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Add116_2_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Add116_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add116_2_impl_out,
                 X => Delay1No126_out_to_Add116_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Add116_2_impl_parent_implementedSystem_port_1_cast);

SharedReg324_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg324_out;
SharedReg265_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg265_out;
SharedReg337_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg337_out;
SharedReg6_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg232_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg232_out;
SharedReg409_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg409_out;
   MUX_Add116_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg324_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg265_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg337_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg232_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Add116_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add116_2_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_2_impl_0_out,
                 Y => Delay1No126_out);

SharedReg726_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg726_out;
SharedReg170_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg170_out;
SharedReg342_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg22_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg531_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg531_out;
SharedReg839_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg839_out;
   MUX_Add116_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg726_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg342_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg531_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg839_out_to_MUX_Add116_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add116_2_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add116_2_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Add117_0_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Add117_0_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Add117_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_0_impl_out,
                 X => Delay1No128_out_to_Add117_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Add117_0_impl_parent_implementedSystem_port_1_cast);

SharedReg368_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg368_out;
SharedReg8_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg259_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg259_out;
SharedReg600_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg600_out;
SharedReg171_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg171_out;
SharedReg302_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg302_out;
   MUX_Add117_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg368_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg259_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg600_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg171_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg302_out_to_MUX_Add117_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_0_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_0_impl_0_out,
                 Y => Delay1No128_out);

SharedReg373_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg373_out;
SharedReg24_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg87_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg87_out;
SharedReg831_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg831_out;
SharedReg274_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg274_out;
SharedReg311_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg311_out;
   MUX_Add117_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg373_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg87_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg831_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg274_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg311_out_to_MUX_Add117_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_0_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_0_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Add117_1_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Add117_1_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Add117_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_1_impl_out,
                 X => Delay1No130_out_to_Add117_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Add117_1_impl_parent_implementedSystem_port_1_cast);

SharedReg304_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg304_out;
SharedReg369_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg369_out;
SharedReg8_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg262_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg149_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg149_out;
SharedReg355_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg355_out;
   MUX_Add117_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg304_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg369_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg8_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg262_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg149_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg355_out_to_MUX_Add117_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_1_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_1_impl_0_out,
                 Y => Delay1No130_out);

SharedReg312_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg312_out;
SharedReg374_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg374_out;
SharedReg24_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg91_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg91_out;
SharedReg152_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg152_out;
SharedReg742_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg742_out;
   MUX_Add117_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg312_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg374_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg91_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg742_out_to_MUX_Add117_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_1_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_1_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Add117_2_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Add117_2_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Add117_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_2_impl_out,
                 X => Delay1No132_out_to_Add117_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Add117_2_impl_parent_implementedSystem_port_1_cast);

SharedReg195_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg195_out;
SharedReg746_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg746_out;
Delay4No57_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_3_cast <= Delay4No57_out;
SharedReg7_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg7_out;
SharedReg251_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg251_out;
SharedReg531_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg531_out;
   MUX_Add117_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg195_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg746_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No57_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg7_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg251_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg531_out_to_MUX_Add117_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_2_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_2_impl_0_out,
                 Y => Delay1No132_out);

SharedReg281_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg281_out;
SharedReg729_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg729_out;
Delay4No62_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No62_out;
SharedReg23_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
SharedReg154_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg157_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg157_out;
   MUX_Add117_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg281_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg729_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No62_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg23_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg157_out_to_MUX_Add117_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_2_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_2_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Add117_3_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Add117_3_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Add117_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add117_3_impl_out,
                 X => Delay1No134_out_to_Add117_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Add117_3_impl_parent_implementedSystem_port_1_cast);

SharedReg412_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg412_out;
SharedReg328_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg328_out;
SharedReg284_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg284_out;
SharedReg338_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg338_out;
SharedReg7_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg253_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg253_out;
   MUX_Add117_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg412_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg328_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg284_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg338_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg253_out_to_MUX_Add117_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_3_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_3_impl_0_out,
                 Y => Delay1No134_out);

SharedReg842_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg842_out;
SharedReg749_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg749_out;
SharedReg181_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg181_out;
SharedReg343_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg23_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg543_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg543_out;
   MUX_Add117_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg842_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg749_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg181_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg543_out_to_MUX_Add117_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add117_3_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add117_3_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Add29_3_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Add29_3_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Add29_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add29_3_impl_out,
                 X => Delay1No136_out_to_Add29_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Add29_3_impl_parent_implementedSystem_port_1_cast);

SharedReg543_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg543_out;
SharedReg205_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg805_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg805_out;
Delay4No58_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_4_cast <= Delay4No58_out;
SharedReg8_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg308_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg308_out;
   MUX_Add29_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg543_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg805_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No58_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg308_out_to_MUX_Add29_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add29_3_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add29_3_impl_0_out,
                 Y => Delay1No136_out);

SharedReg48_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg534_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg534_out;
SharedReg753_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg753_out;
Delay4No63_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_4_cast <= Delay4No63_out;
SharedReg24_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg297_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg297_out;
   MUX_Add29_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg534_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg753_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No63_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg297_out_to_MUX_Add29_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add29_3_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add29_3_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Add36_4_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Add36_4_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Add36_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add36_4_impl_out,
                 X => Delay1No138_out_to_Add36_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Add36_4_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg310_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg310_out;
SharedReg596_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg596_out;
SharedReg332_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg332_out;
SharedReg310_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg310_out;
Delay4No79_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_6_cast <= Delay4No79_out;
   MUX_Add36_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg310_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg596_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg332_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg310_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No79_out_to_MUX_Add36_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add36_4_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add36_4_impl_0_out,
                 Y => Delay1No138_out);

SharedReg25_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg299_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg299_out;
SharedReg846_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg846_out;
SharedReg734_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg734_out;
SharedReg315_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg315_out;
Delay4No84_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No84_out;
   MUX_Add36_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg299_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg846_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg734_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg315_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No84_out_to_MUX_Add36_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add36_4_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add36_4_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Add126_0_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Add126_0_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Add126_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add126_0_impl_out,
                 X => Delay1No140_out_to_Add126_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Add126_0_impl_parent_implementedSystem_port_1_cast);

Delay4No75_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No75_out;
SharedReg9_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg302_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg302_out;
SharedReg87_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg87_out;
SharedReg351_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg340_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg340_out;
   MUX_Add126_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No75_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg302_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg87_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg340_out_to_MUX_Add126_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add126_0_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add126_0_impl_0_out,
                 Y => Delay1No140_out);

Delay4No80_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No80_out;
SharedReg25_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg291_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg291_out;
SharedReg541_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg541_out;
SharedReg738_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg738_out;
SharedReg345_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg345_out;
   MUX_Add126_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No80_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg291_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg541_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg738_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg345_out_to_MUX_Add126_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add126_0_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add126_0_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Add126_4_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Add126_4_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Add126_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add126_4_impl_out,
                 X => Delay1No142_out_to_Add126_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Add126_4_impl_parent_implementedSystem_port_1_cast);

SharedReg10_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg372_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg827_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg827_out;
SharedReg185_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg185_out;
SharedReg344_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg344_out;
SharedReg432_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg432_out;
   MUX_Add126_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg827_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg185_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg344_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg432_out_to_MUX_Add126_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add126_4_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add126_4_impl_0_out,
                 Y => Delay1No142_out);

SharedReg26_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg377_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg377_out;
SharedReg549_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg549_out;
SharedReg476_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg476_out;
SharedReg349_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg349_out;
SharedReg461_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg461_out;
   MUX_Add126_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg377_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg549_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg476_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg349_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg461_out_to_MUX_Add126_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add126_4_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add126_4_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Add37_2_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Add37_2_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Add37_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add37_2_impl_out,
                 X => Delay1No144_out_to_Add37_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Add37_2_impl_parent_implementedSystem_port_1_cast);

SharedReg358_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg358_out;
SharedReg306_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg306_out;
SharedReg370_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg370_out;
SharedReg8_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg8_out;
SharedReg306_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg306_out;
Delay2No322_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_6_cast <= Delay2No322_out;
   MUX_Add37_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg358_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg306_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg370_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg8_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg306_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay2No322_out_to_MUX_Add37_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add37_2_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add37_2_impl_0_out,
                 Y => Delay1No144_out);

SharedReg803_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg313_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg313_out;
SharedReg375_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg375_out;
SharedReg24_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg24_out;
SharedReg295_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg295_out;
Delay2No327_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_6_cast <= Delay2No327_out;
   MUX_Add37_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg313_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg375_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg24_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg295_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay2No327_out_to_MUX_Add37_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add37_2_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add37_2_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Add127_1_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Add127_1_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Add127_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_1_impl_out,
                 X => Delay1No146_out_to_Add127_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Add127_1_impl_parent_implementedSystem_port_1_cast);

SharedReg341_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg341_out;
Delay4No76_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No76_out;
SharedReg9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg304_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg304_out;
Delay2No321_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_5_cast <= Delay2No321_out;
SharedReg214_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg214_out;
   MUX_Add127_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg341_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No76_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg304_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay2No321_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg214_out_to_MUX_Add127_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add127_1_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_1_impl_0_out,
                 Y => Delay1No146_out);

SharedReg346_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg346_out;
Delay4No81_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No81_out;
SharedReg25_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg293_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg293_out;
Delay2No326_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_5_cast <= Delay2No326_out;
SharedReg526_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg526_out;
   MUX_Add127_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No81_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg25_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg293_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay2No326_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg526_out_to_MUX_Add127_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add127_1_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_1_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Add127_2_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Add127_2_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Add127_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_2_impl_out,
                 X => Delay1No148_out_to_Add127_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Add127_2_impl_parent_implementedSystem_port_1_cast);

SharedReg218_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg218_out;
SharedReg342_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg342_out;
Delay4No77_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_3_cast <= Delay4No77_out;
SharedReg9_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg9_out;
SharedReg370_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg370_out;
SharedReg337_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg337_out;
   MUX_Add127_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg218_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg342_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No77_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg9_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg370_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg337_out_to_MUX_Add127_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add127_2_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_2_impl_0_out,
                 Y => Delay1No148_out);

SharedReg530_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg530_out;
SharedReg347_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg347_out;
Delay4No82_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No82_out;
SharedReg25_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg375_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg375_out;
SharedReg305_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg305_out;
   MUX_Add127_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg530_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg347_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No82_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg375_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg305_out_to_MUX_Add127_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add127_2_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_2_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Add127_3_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Add127_3_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Add127_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_3_impl_out,
                 X => Delay1No150_out_to_Add127_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Add127_3_impl_parent_implementedSystem_port_1_cast);

Delay2No323_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_1_cast <= Delay2No323_out;
SharedReg361_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg361_out;
SharedReg308_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg308_out;
SharedReg371_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg371_out;
SharedReg9_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg9_out;
SharedReg371_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg371_out;
   MUX_Add127_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No323_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg361_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg308_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg371_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg9_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg371_out_to_MUX_Add127_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add127_3_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_3_impl_0_out,
                 Y => Delay1No150_out);

Delay2No328_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_1_cast <= Delay2No328_out;
SharedReg847_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg847_out;
SharedReg314_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg314_out;
SharedReg376_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg376_out;
SharedReg25_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg25_out;
SharedReg376_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg376_out;
   MUX_Add127_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No328_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg847_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg314_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg376_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg25_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg376_out_to_MUX_Add127_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add127_3_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_3_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Add38_0_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Add38_0_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Add38_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add38_0_impl_out,
                 X => Delay1No152_out_to_Add38_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Add38_0_impl_parent_implementedSystem_port_1_cast);

SharedReg424_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg424_out;
SharedReg10_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg368_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg368_out;
Delay2No320_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_4_cast <= Delay2No320_out;
SharedReg224_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg368_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg368_out;
   MUX_Add38_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg424_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg368_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No320_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg368_out_to_MUX_Add38_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_0_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_0_impl_0_out,
                 Y => Delay1No152_out);

SharedReg453_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg453_out;
SharedReg26_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg373_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg373_out;
Delay2No325_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_4_cast <= Delay2No325_out;
SharedReg522_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg522_out;
SharedReg373_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg373_out;
   MUX_Add38_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg453_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg373_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No325_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg522_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg373_out_to_MUX_Add38_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_0_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_0_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Add38_1_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Add38_1_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Add38_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add38_1_impl_out,
                 X => Delay1No154_out_to_Add38_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Add38_1_impl_parent_implementedSystem_port_1_cast);

SharedReg369_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg369_out;
SharedReg426_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg426_out;
SharedReg10_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg10_out;
SharedReg369_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg369_out;
SharedReg336_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg336_out;
SharedReg336_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg336_out;
   MUX_Add38_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg369_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg426_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg10_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg369_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg336_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg336_out_to_MUX_Add38_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_1_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_1_impl_0_out,
                 Y => Delay1No154_out);

SharedReg374_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg374_out;
SharedReg455_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg455_out;
SharedReg26_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg374_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg374_out;
SharedReg303_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg303_out;
SharedReg341_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg341_out;
   MUX_Add38_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg374_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg455_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg26_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg374_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg303_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg341_out_to_MUX_Add38_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_1_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_1_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Add38_2_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Add38_2_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Add38_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add38_2_impl_out,
                 X => Delay1No156_out_to_Add38_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Add38_2_impl_parent_implementedSystem_port_1_cast);

SharedReg337_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg337_out;
SharedReg370_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg370_out;
SharedReg428_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg428_out;
SharedReg10_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg429_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg429_out;
SharedReg578_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg578_out;
   MUX_Add38_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg337_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg370_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg428_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg10_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg429_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg578_out_to_MUX_Add38_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_2_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_2_impl_0_out,
                 Y => Delay1No156_out);

SharedReg342_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg342_out;
SharedReg375_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg375_out;
SharedReg457_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg457_out;
SharedReg26_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg458_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg458_out;
SharedReg515_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg515_out;
   MUX_Add38_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg342_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg375_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg457_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg458_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg515_out_to_MUX_Add38_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_2_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_2_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Add38_3_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Add38_3_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Add38_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add38_3_impl_out,
                 X => Delay1No158_out_to_Add38_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Add38_3_impl_parent_implementedSystem_port_1_cast);

SharedReg338_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg338_out;
SharedReg237_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg237_out;
SharedReg343_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg343_out;
Delay4No78_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_4_cast <= Delay4No78_out;
SharedReg10_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg10_out;
SharedReg431_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg431_out;
   MUX_Add38_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg338_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg237_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg343_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No78_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg10_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg431_out_to_MUX_Add38_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_3_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_3_impl_0_out,
                 Y => Delay1No158_out);

SharedReg307_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg307_out;
SharedReg542_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg542_out;
SharedReg348_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg348_out;
Delay4No83_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_4_cast <= Delay4No83_out;
SharedReg26_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg26_out;
SharedReg460_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg460_out;
   MUX_Add38_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg307_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg542_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg348_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No83_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg26_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg460_out_to_MUX_Add38_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add38_3_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add38_3_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Add128_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_0_impl_out,
                 X => Delay1No160_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast);

SharedReg490_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg490_out;
SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
SharedReg425_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg425_out;
SharedReg335_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg335_out;
SharedReg335_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg335_out;
SharedReg414_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg414_out;
   MUX_Add128_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg490_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg425_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg335_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg335_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg414_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_0_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_0_impl_0_out,
                 Y => Delay1No160_out);

SharedReg500_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg500_out;
SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg454_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg454_out;
SharedReg301_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg301_out;
SharedReg340_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg340_out;
SharedReg425_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg425_out;
   MUX_Add128_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg500_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg454_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg301_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg340_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg425_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_0_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_0_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Add128_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_1_impl_out,
                 X => Delay1No162_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast);

SharedReg416_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg416_out;
SharedReg492_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg492_out;
SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg427_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg427_out;
SharedReg575_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg575_out;
SharedReg369_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg369_out;
   MUX_Add128_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg416_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg492_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg427_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg575_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg369_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_1_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_1_impl_0_out,
                 Y => Delay1No162_out);

SharedReg427_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg502_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg502_out;
SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg456_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg456_out;
SharedReg513_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg513_out;
SharedReg374_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg374_out;
   MUX_Add128_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg502_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg456_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg513_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg374_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_1_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_1_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Add128_2_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Add128_2_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Add128_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_2_impl_out,
                 X => Delay1No164_out_to_Add128_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Add128_2_impl_parent_implementedSystem_port_1_cast);

SharedReg370_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg370_out;
SharedReg418_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg418_out;
SharedReg494_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg494_out;
SharedReg11_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg428_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg428_out;
SharedReg555_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg555_out;
   MUX_Add128_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg370_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg418_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg494_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg428_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg555_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_2_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_2_impl_0_out,
                 Y => Delay1No164_out);

SharedReg375_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg375_out;
SharedReg429_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg504_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg504_out;
SharedReg27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg27_out;
SharedReg457_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg457_out;
SharedReg347_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg347_out;
   MUX_Add128_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg375_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg504_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg457_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg347_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_2_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_2_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Add128_3_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Add128_3_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Add128_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_3_impl_out,
                 X => Delay1No166_out_to_Add128_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Add128_3_impl_parent_implementedSystem_port_1_cast);

SharedReg581_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg581_out;
SharedReg338_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg371_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg371_out;
SharedReg430_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg430_out;
SharedReg11_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg11_out;
SharedReg430_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg430_out;
   MUX_Add128_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg581_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg371_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg430_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg11_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg430_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_3_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_3_impl_0_out,
                 Y => Delay1No166_out);

SharedReg517_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg517_out;
SharedReg343_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg343_out;
SharedReg376_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg376_out;
SharedReg459_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg459_out;
SharedReg27_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg27_out;
SharedReg459_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg459_out;
   MUX_Add128_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg517_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg343_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg376_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg459_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg27_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg459_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_3_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_3_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Add128_4_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Add128_4_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Add128_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_4_impl_out,
                 X => Delay1No168_out_to_Add128_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Add128_4_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg433_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg433_out;
Delay2No324_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_3_cast <= Delay2No324_out;
SharedReg333_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg333_out;
SharedReg372_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg372_out;
SharedReg498_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg498_out;
   MUX_Add128_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg433_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No324_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg333_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg372_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg498_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_4_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_4_impl_0_out,
                 Y => Delay1No168_out);

SharedReg27_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg462_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg462_out;
Delay2No329_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_3_cast <= Delay2No329_out;
SharedReg808_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg377_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg377_out;
SharedReg508_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg508_out;
   MUX_Add128_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg462_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No329_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg377_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg508_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add128_4_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_4_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Add129_0_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Add129_0_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Add129_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_0_impl_out,
                 X => Delay1No170_out_to_Add129_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Add129_0_impl_parent_implementedSystem_port_1_cast);

Delay4No90_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No90_out;
SharedReg13_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg424_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg424_out;
SharedReg572_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg572_out;
SharedReg368_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg368_out;
SharedReg463_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg463_out;
   MUX_Add129_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No90_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg424_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg572_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg368_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg463_out_to_MUX_Add129_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_0_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_0_impl_0_out,
                 Y => Delay1No170_out);

Delay4No95_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No95_out;
SharedReg29_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg453_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg453_out;
SharedReg511_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg511_out;
SharedReg373_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg373_out;
SharedReg480_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg480_out;
   MUX_Add129_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No95_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg453_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg511_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg373_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg480_out_to_MUX_Add129_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_0_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_0_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Add129_1_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Add129_1_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Add129_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_1_impl_out,
                 X => Delay1No172_out_to_Add129_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Add129_1_impl_parent_implementedSystem_port_1_cast);

SharedReg465_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg465_out;
Delay4No91_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No91_out;
SharedReg13_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg426_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg426_out;
SharedReg553_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg553_out;
SharedReg492_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg492_out;
   MUX_Add129_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg465_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No91_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg13_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg426_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg553_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg492_out_to_MUX_Add129_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_1_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_1_impl_0_out,
                 Y => Delay1No172_out);

SharedReg482_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg482_out;
Delay4No96_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No96_out;
SharedReg29_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg455_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg455_out;
SharedReg346_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg346_out;
SharedReg502_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg502_out;
   MUX_Add129_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg482_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No96_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg29_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg455_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg346_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg502_out_to_MUX_Add129_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_1_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_1_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Add129_2_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Add129_2_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Add129_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_2_impl_out,
                 X => Delay1No174_out_to_Add129_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Add129_2_impl_parent_implementedSystem_port_1_cast);

SharedReg494_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg494_out;
SharedReg467_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg467_out;
Delay4No92_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_3_cast <= Delay4No92_out;
SharedReg13_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg13_out;
SharedReg495_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg495_out;
SharedReg667_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg667_out;
   MUX_Add129_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg494_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg467_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No92_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg13_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg495_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg667_out_to_MUX_Add129_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_2_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_2_impl_0_out,
                 Y => Delay1No174_out);

SharedReg504_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg484_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg484_out;
Delay4No97_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No97_out;
SharedReg29_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg29_out;
SharedReg505_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg505_out;
SharedReg711_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg711_out;
   MUX_Add129_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg484_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No97_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg29_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg505_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg711_out_to_MUX_Add129_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_2_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_2_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Add129_3_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Add129_3_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Add129_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_3_impl_out,
                 X => Delay1No176_out_to_Add129_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Add129_3_impl_parent_implementedSystem_port_1_cast);

SharedReg557_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg557_out;
SharedReg371_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg371_out;
SharedReg420_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg420_out;
SharedReg496_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg496_out;
SharedReg13_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg497_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg497_out;
   MUX_Add129_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg557_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg371_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg420_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg496_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg497_out_to_MUX_Add129_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_3_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_3_impl_0_out,
                 Y => Delay1No176_out);

SharedReg348_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg376_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg376_out;
SharedReg431_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg431_out;
SharedReg506_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg506_out;
SharedReg29_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg29_out;
SharedReg507_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg507_out;
   MUX_Add129_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg376_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg431_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg506_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg29_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg507_out_to_MUX_Add129_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_3_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_3_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Add129_4_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Add129_4_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Add129_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_4_impl_out,
                 X => Delay1No178_out_to_Add129_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Add129_4_impl_parent_implementedSystem_port_1_cast);

SharedReg13_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg432_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg432_out;
SharedReg339_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg339_out;
SharedReg271_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg271_out;
SharedReg422_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg422_out;
Delay4No94_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_6_cast <= Delay4No94_out;
   MUX_Add129_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg432_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg339_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg271_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg422_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No94_out_to_MUX_Add129_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_4_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_4_impl_0_out,
                 Y => Delay1No178_out);

SharedReg29_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg29_out;
SharedReg461_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg461_out;
SharedReg309_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg309_out;
SharedReg546_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg546_out;
SharedReg433_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg433_out;
Delay4No99_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No99_out;
   MUX_Add129_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg461_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg309_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg546_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg433_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No99_out_to_MUX_Add129_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add129_4_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_4_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Add40_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_0_impl_out,
                 X => Delay1No180_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast);

SharedReg560_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg560_out;
SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg491_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg491_out;
SharedReg551_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg551_out;
SharedReg490_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg490_out;
Delay3No200_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast <= Delay3No200_out;
   MUX_Add40_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg560_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg491_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg551_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg490_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No200_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_0_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_0_impl_0_out,
                 Y => Delay1No180_out);

SharedReg570_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg570_out;
SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg501_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg501_out;
SharedReg345_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg345_out;
SharedReg500_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg500_out;
Delay3No205_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast <= Delay3No205_out;
   MUX_Add40_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg570_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg501_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg345_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg500_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No205_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_0_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_0_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Add40_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_1_impl_out,
                 X => Delay1No182_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast);

Delay3No201_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No201_out;
SharedReg562_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg493_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg493_out;
SharedReg665_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg665_out;
SharedReg562_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg562_out;
   MUX_Add40_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No201_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg493_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg665_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg562_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_1_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_1_impl_0_out,
                 Y => Delay1No182_out);

Delay3No206_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast <= Delay3No206_out;
SharedReg573_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg573_out;
SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg503_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg503_out;
SharedReg709_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg709_out;
SharedReg573_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg573_out;
   MUX_Add40_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No206_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg573_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg503_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg709_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg573_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_1_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_1_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Add40_2_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Add40_2_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Add40_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_2_impl_out,
                 X => Delay1No184_out_to_Add40_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Add40_2_impl_parent_implementedSystem_port_1_cast);

SharedReg564_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg564_out;
Delay3No202_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_2_cast <= Delay3No202_out;
SharedReg564_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg564_out;
SharedReg14_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg555_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg555_out;
SharedReg762_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg762_out;
   MUX_Add40_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg564_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No202_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg564_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg14_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg555_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg762_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_2_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_2_impl_0_out,
                 Y => Delay1No184_out);

SharedReg576_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg576_out;
Delay3No207_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_2_cast <= Delay3No207_out;
SharedReg576_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg576_out;
SharedReg30_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg30_out;
SharedReg494_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg494_out;
SharedReg773_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg773_out;
   MUX_Add40_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg576_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No207_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg576_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg30_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg494_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg773_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_2_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_2_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Add40_3_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Add40_3_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Add40_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_3_impl_out,
                 X => Delay1No186_out_to_Add40_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Add40_3_impl_parent_implementedSystem_port_1_cast);

SharedReg669_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg669_out;
SharedReg496_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg496_out;
SharedReg469_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg469_out;
Delay4No93_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_4_cast <= Delay4No93_out;
SharedReg14_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg14_out;
SharedReg557_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg557_out;
   MUX_Add40_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg669_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg496_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg469_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No93_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg14_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg557_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_3_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_3_impl_0_out,
                 Y => Delay1No186_out);

SharedReg713_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg713_out;
SharedReg506_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg506_out;
SharedReg486_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg486_out;
Delay4No98_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_4_cast <= Delay4No98_out;
SharedReg30_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg496_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg496_out;
   MUX_Add40_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg713_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg506_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg486_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No98_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg496_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_3_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_3_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Add40_4_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Add40_4_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Add40_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_4_impl_out,
                 X => Delay1No188_out_to_Add40_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Add40_4_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg499_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg499_out;
SharedReg584_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg584_out;
SharedReg339_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg339_out;
SharedReg471_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg471_out;
SharedReg568_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg568_out;
   MUX_Add40_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg499_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg584_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg339_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg471_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg568_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_4_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_4_impl_0_out,
                 Y => Delay1No188_out);

SharedReg30_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg30_out;
SharedReg509_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg509_out;
SharedReg519_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg519_out;
SharedReg344_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg344_out;
SharedReg488_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg488_out;
SharedReg582_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg582_out;
   MUX_Add40_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg30_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg509_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg519_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg344_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg488_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg582_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add40_4_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_4_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Add130_0_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Add130_0_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Add130_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_0_impl_out,
                 X => Delay1No190_out_to_Add130_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Add130_0_impl_parent_implementedSystem_port_1_cast);

SharedReg673_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg673_out;
SharedReg15_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg551_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg551_out;
SharedReg663_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg663_out;
SharedReg560_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg560_out;
SharedReg510_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg510_out;
   MUX_Add130_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg673_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg551_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg663_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg560_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg510_out_to_MUX_Add130_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_0_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_0_impl_0_out,
                 Y => Delay1No190_out);

SharedReg683_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg683_out;
SharedReg31_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg490_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg490_out;
SharedReg707_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg707_out;
SharedReg570_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg570_out;
SharedReg550_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg550_out;
   MUX_Add130_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg683_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg490_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg707_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg570_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg550_out_to_MUX_Add130_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_0_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_0_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Add130_1_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Add130_1_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Add130_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_1_impl_out,
                 X => Delay1No192_out_to_Add130_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Add130_1_impl_parent_implementedSystem_port_1_cast);

SharedReg512_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg512_out;
SharedReg675_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg675_out;
SharedReg15_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg15_out;
SharedReg553_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg553_out;
SharedReg760_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg760_out;
SharedReg689_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg689_out;
   MUX_Add130_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg512_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg675_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg15_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg553_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg760_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg689_out_to_MUX_Add130_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_1_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_1_impl_0_out,
                 Y => Delay1No192_out);

SharedReg552_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg552_out;
SharedReg684_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg684_out;
SharedReg31_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg492_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg492_out;
SharedReg771_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg771_out;
SharedReg698_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg698_out;
   MUX_Add130_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg552_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg684_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg31_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg492_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg771_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg698_out_to_MUX_Add130_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_1_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_1_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Add130_2_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Add130_2_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Add130_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_2_impl_out,
                 X => Delay1No194_out_to_Add130_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Add130_2_impl_parent_implementedSystem_port_1_cast);

SharedReg690_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg690_out;
SharedReg514_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg514_out;
SharedReg677_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg677_out;
SharedReg15_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg15_out;
SharedReg701_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg701_out;
SharedReg428_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg428_out;
   MUX_Add130_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg690_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg514_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg677_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg15_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg701_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg428_out_to_MUX_Add130_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_2_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_2_impl_0_out,
                 Y => Delay1No194_out);

SharedReg700_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg700_out;
SharedReg554_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg554_out;
SharedReg685_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg685_out;
SharedReg31_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg31_out;
SharedReg589_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg589_out;
SharedReg457_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg457_out;
   MUX_Add130_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg700_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg554_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg685_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg31_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg589_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg457_out_to_MUX_Add130_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_2_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_2_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Add130_3_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Add130_3_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Add130_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_3_impl_out,
                 X => Delay1No196_out_to_Add130_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Add130_3_impl_parent_implementedSystem_port_1_cast);

SharedReg764_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg764_out;
SharedReg566_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg566_out;
Delay3No203_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_3_cast <= Delay3No203_out;
SharedReg566_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg566_out;
SharedReg15_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg703_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg703_out;
   MUX_Add130_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg764_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg566_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No203_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg566_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg15_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg703_out_to_MUX_Add130_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_3_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_3_impl_0_out,
                 Y => Delay1No196_out);

SharedReg775_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg775_out;
SharedReg579_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg579_out;
Delay3No208_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_3_cast <= Delay3No208_out;
SharedReg579_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg579_out;
SharedReg31_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg31_out;
SharedReg591_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg591_out;
   MUX_Add130_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg775_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg579_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No208_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg579_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg31_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg591_out_to_MUX_Add130_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_3_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_3_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Add130_4_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Add130_4_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Add130_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_4_impl_out,
                 X => Delay1No198_out_to_Add130_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Add130_4_impl_parent_implementedSystem_port_1_cast);

SharedReg15_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg559_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg559_out;
SharedReg559_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg559_out;
SharedReg372_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg372_out;
Delay3No204_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_5_cast <= Delay3No204_out;
SharedReg681_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg681_out;
   MUX_Add130_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg559_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg559_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg372_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No204_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg681_out_to_MUX_Add130_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_4_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_4_impl_0_out,
                 Y => Delay1No198_out);

SharedReg31_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg31_out;
SharedReg498_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg498_out;
SharedReg349_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg349_out;
SharedReg377_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg377_out;
Delay3No209_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_5_cast <= Delay3No209_out;
SharedReg687_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg687_out;
   MUX_Add130_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg31_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg498_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg349_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg377_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No209_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg687_out_to_MUX_Add130_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add130_4_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_4_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No200_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg49_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg900_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg944_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg944_out;
SharedReg171_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg171_out;
SharedReg913_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg64_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg64_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg944_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg171_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg64_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No200_out);

SharedReg909_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg830_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg830_out;
SharedReg912_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg162_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg162_out;
SharedReg914_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg914_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg830_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg162_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg914_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No202_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg67_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg67_out;
SharedReg52_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg52_out;
SharedReg900_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg944_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg944_out;
SharedReg164_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg164_out;
SharedReg913_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg67_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg52_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg944_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg164_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No202_out);

SharedReg914_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg914_out;
SharedReg909_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg834_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg834_out;
SharedReg912_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg159_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg159_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg914_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg834_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg159_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No204_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg69_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg55_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg900_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg944_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg944_out;
SharedReg177_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg177_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg944_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg177_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No204_out);

SharedReg168_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg168_out;
SharedReg914_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg914_out;
SharedReg909_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg39_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg39_out;
SharedReg838_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg838_out;
SharedReg912_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg168_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg914_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg39_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg838_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No206_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg182_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg913_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg82_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg57_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg57_out;
SharedReg900_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg944_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg944_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg82_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg57_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg944_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No206_out);

SharedReg912_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg180_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg180_out;
SharedReg914_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg914_out;
SharedReg909_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg42_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg42_out;
SharedReg822_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg822_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg180_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg914_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg42_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg822_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No208_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg944_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg944_out;
SharedReg191_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg191_out;
SharedReg913_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg84_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg84_out;
SharedReg60_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg60_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg944_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg191_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg84_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg60_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No208_out);

SharedReg46_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg845_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg845_out;
SharedReg912_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg186_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg186_out;
SharedReg914_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg914_out;
SharedReg909_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg845_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg186_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg914_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product11_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_0_impl_out,
                 X => Delay1No210_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg799_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg940_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg940_out;
SharedReg902_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg914_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg914_out;
   MUX_Product11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg940_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg914_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_0_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_0_impl_0_out,
                 Y => Delay1No210_out);

SharedReg49_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg924_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg924_out;
SharedReg830_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg830_out;
SharedReg171_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg171_out;
SharedReg162_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg162_out;
SharedReg50_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg50_out;
   MUX_Product11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg924_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg830_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg171_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg162_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg50_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_0_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_0_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product11_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_1_impl_out,
                 X => Delay1No212_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg914_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg914_out;
SharedReg899_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg802_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg802_out;
SharedReg940_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg940_out;
SharedReg902_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg914_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg802_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg940_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_1_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_0_out,
                 Y => Delay1No212_out);

SharedReg53_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg52_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg52_out;
SharedReg924_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg924_out;
SharedReg834_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg834_out;
SharedReg164_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg164_out;
SharedReg159_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg159_out;
   MUX_Product11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg52_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg924_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg834_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg164_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg159_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_1_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product11_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_2_impl_out,
                 X => Delay1No214_out_to_Product11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg914_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg914_out;
SharedReg899_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg859_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg859_out;
SharedReg940_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg940_out;
SharedReg902_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg914_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg859_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg940_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_2_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_2_impl_0_out,
                 Y => Delay1No214_out);

SharedReg168_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg168_out;
SharedReg56_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg56_out;
SharedReg55_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg924_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg924_out;
SharedReg838_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg838_out;
SharedReg177_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg177_out;
   MUX_Product11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg168_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg56_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg924_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg838_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg177_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_2_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_2_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Product11_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_3_impl_out,
                 X => Delay1No216_out_to_Product11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Product11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg914_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg914_out;
SharedReg899_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg848_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg848_out;
SharedReg940_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg940_out;
   MUX_Product11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg914_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg848_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg940_out_to_MUX_Product11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_3_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_3_impl_0_out,
                 Y => Delay1No216_out);

SharedReg182_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg180_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg180_out;
SharedReg71_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg71_out;
SharedReg57_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg57_out;
SharedReg924_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg924_out;
SharedReg822_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg822_out;
   MUX_Product11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg180_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg71_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg57_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg924_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg822_out_to_MUX_Product11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_3_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_3_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Product11_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_4_impl_out,
                 X => Delay1No218_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg809_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg809_out;
SharedReg940_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg940_out;
SharedReg902_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg914_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg914_out;
SharedReg899_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg809_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg940_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg914_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_4_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_0_out,
                 Y => Delay1No218_out);

SharedReg924_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg924_out;
SharedReg845_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg845_out;
SharedReg191_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg191_out;
SharedReg186_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg186_out;
SharedReg73_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg73_out;
SharedReg60_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg60_out;
   MUX_Product11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg924_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg845_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg191_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg186_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg73_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg60_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product11_4_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No220_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg904_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg904_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No220_out);

SharedReg63_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg50_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg50_out;
SharedReg188_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg188_out;
SharedReg64_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg64_out;
SharedReg50_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg50_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg50_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg188_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg50_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product21_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_1_impl_out,
                 X => Delay1No222_out_to_Product21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg904_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg904_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_1_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_0_out,
                 Y => Delay1No222_out);

SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg66_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg36_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg174_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg174_out;
SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg53_out;
   MUX_Product21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg174_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg53_out_to_MUX_Product21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_1_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_1_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product21_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_2_impl_out,
                 X => Delay1No224_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg904_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_2_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_0_out,
                 Y => Delay1No224_out);

SharedReg56_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg56_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg56_out;
SharedReg68_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg39_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg39_out;
SharedReg39_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg195_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg195_out;
   MUX_Product21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg56_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg39_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_2_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Product21_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_3_impl_out,
                 X => Delay1No226_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg904_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_3_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_0_out,
                 Y => Delay1No226_out);

SharedReg205_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg205_out;
SharedReg71_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg71_out;
SharedReg71_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg71_out;
SharedReg70_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg70_out;
SharedReg42_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg42_out;
SharedReg42_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg42_out;
   MUX_Product21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg205_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg71_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg70_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg42_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg42_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_3_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Product21_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_4_impl_out,
                 X => Delay1No228_out_to_Product21_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Product21_4_impl_parent_implementedSystem_port_1_cast);

SharedReg910_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product21_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg904_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product21_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_4_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_0_out,
                 Y => Delay1No228_out);

SharedReg46_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg241_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg241_out;
SharedReg95_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg73_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg73_out;
SharedReg72_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg72_out;
   MUX_Product21_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg241_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg73_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg72_out_to_MUX_Product21_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product21_4_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_4_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No230_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg311_out;
SharedReg363_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg363_out;
SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg311_out;
SharedReg697_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg697_out;
SharedReg363_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg363_out;
SharedReg291_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg291_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg363_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg311_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg697_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg363_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg291_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No230_out);

SharedReg345_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg345_out;
SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg378_out;
SharedReg345_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg673_out;
SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg378_out;
SharedReg292_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg292_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg345_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg345_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg673_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg378_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg292_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No232_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg293_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg293_out;
SharedReg312_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg312_out;
SharedReg364_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg364_out;
SharedReg312_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg312_out;
SharedReg761_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg761_out;
SharedReg482_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg482_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg293_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg364_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg312_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg761_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg482_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No232_out);

SharedReg294_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg294_out;
SharedReg346_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg379_out;
SharedReg346_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg346_out;
SharedReg770_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg770_out;
SharedReg512_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg512_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg294_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg346_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg770_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg512_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No234_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg484_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg484_out;
SharedReg295_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg295_out;
SharedReg313_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg313_out;
SharedReg365_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg365_out;
SharedReg365_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg365_out;
SharedReg418_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg418_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg484_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg295_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg313_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg365_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg365_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg418_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No234_out);

SharedReg514_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg514_out;
SharedReg296_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg296_out;
SharedReg347_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg347_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg380_out;
SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg467_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg467_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg514_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg296_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg347_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg380_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg467_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No236_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg420_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg420_out;
SharedReg486_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg486_out;
SharedReg297_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg297_out;
SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg314_out;
SharedReg669_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg669_out;
SharedReg421_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg421_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg420_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg486_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg297_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg669_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg421_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No236_out);

SharedReg469_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg469_out;
SharedReg516_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg516_out;
SharedReg298_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg298_out;
SharedReg348_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg348_out;
SharedReg691_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg691_out;
SharedReg470_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg470_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg469_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg516_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg298_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg348_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg691_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg470_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No238_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg671_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg671_out;
SharedReg367_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg367_out;
SharedReg705_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg705_out;
SharedReg315_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg315_out;
SharedReg299_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg299_out;
Delay4No54_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= Delay4No54_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg671_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg367_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg705_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg315_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg299_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No54_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No238_out);

SharedReg692_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg692_out;
SharedReg382_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg382_out;
SharedReg681_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg681_out;
SharedReg349_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg349_out;
SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg300_out;
Delay4No69_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No69_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg692_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg382_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg681_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No69_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Product12_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_0_impl_out,
                 X => Delay1No240_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg923_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg923_out;
SharedReg906_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg904_out;
   MUX_Product12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg923_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg904_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_0_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_0_out,
                 Y => Delay1No240_out);

SharedReg75_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg739_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg739_out;
SharedReg64_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg64_out;
SharedReg209_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg76_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg76_out;
SharedReg64_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg64_out;
   MUX_Product12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg739_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg64_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg76_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg64_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_0_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Product12_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_1_impl_out,
                 X => Delay1No242_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg904_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg923_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg923_out;
SharedReg906_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg904_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg923_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_1_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_0_out,
                 Y => Delay1No242_out);

SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg67_out;
SharedReg77_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg743_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg743_out;
SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg67_out;
SharedReg199_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg199_out;
SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg67_out;
   MUX_Product12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg743_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg199_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_1_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Product12_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_2_impl_out,
                 X => Delay1No244_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg923_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg923_out;
SharedReg906_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg904_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg923_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_2_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_0_out,
                 Y => Delay1No244_out);

SharedReg69_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg69_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg79_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg804_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg804_out;
SharedReg56_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg56_out;
SharedReg202_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg202_out;
   MUX_Product12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg79_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg804_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg56_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg202_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_2_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product12_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_3_impl_out,
                 X => Delay1No246_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg923_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg923_out;
SharedReg906_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg904_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg923_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_3_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_0_out,
                 Y => Delay1No246_out);

SharedReg221_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg82_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg82_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg81_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg81_out;
SharedReg805_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg805_out;
SharedReg58_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg58_out;
   MUX_Product12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg82_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg81_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg805_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg58_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_3_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Product12_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_4_impl_out,
                 X => Delay1No248_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg923_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg923_out;
SharedReg906_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg904_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg904_out;
SharedReg899_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg923_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg904_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_4_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_0_out,
                 Y => Delay1No248_out);

SharedReg755_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg755_out;
SharedReg73_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg73_out;
SharedReg257_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg257_out;
SharedReg97_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg97_out;
SharedReg84_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg84_out;
SharedReg83_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg83_out;
   MUX_Product12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg755_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg257_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg97_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg84_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg83_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product12_4_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Product22_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_0_impl_out,
                 X => Delay1No250_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast);

SharedReg909_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg923_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg923_out;
SharedReg916_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg927_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg927_out;
   MUX_Product22_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg923_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg927_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_0_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_0_impl_0_out,
                 Y => Delay1No250_out);

SharedReg63_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg799_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg50_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg50_out;
SharedReg188_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg188_out;
SharedReg64_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg64_out;
SharedReg866_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg866_out;
   MUX_Product22_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg50_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg188_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg64_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg866_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_0_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_0_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Product22_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_1_impl_out,
                 X => Delay1No252_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast);

SharedReg927_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg927_out;
SharedReg909_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg923_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg923_out;
SharedReg916_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product22_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg927_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg923_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_1_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_1_impl_0_out,
                 Y => Delay1No252_out);

SharedReg868_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg868_out;
SharedReg66_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg802_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg802_out;
SharedReg53_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg53_out;
SharedReg174_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg174_out;
SharedReg53_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg53_out;
   MUX_Product22_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg868_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg802_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg174_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg53_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_1_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_1_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Product22_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_2_impl_out,
                 X => Delay1No254_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg927_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg927_out;
SharedReg909_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg923_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg923_out;
SharedReg916_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product22_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg927_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg923_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_2_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_2_impl_0_out,
                 Y => Delay1No254_out);

SharedReg56_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg870_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg870_out;
SharedReg68_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg859_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg859_out;
SharedReg39_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg39_out;
SharedReg195_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg195_out;
   MUX_Product22_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg870_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg68_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg859_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg39_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg195_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_2_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_2_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Product22_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_3_impl_out,
                 X => Delay1No256_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast);

SharedReg912_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg927_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg927_out;
SharedReg909_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg923_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg923_out;
SharedReg916_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product22_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg927_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg923_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_3_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_3_impl_0_out,
                 Y => Delay1No256_out);

SharedReg205_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg205_out;
SharedReg71_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg71_out;
SharedReg872_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg872_out;
SharedReg70_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg70_out;
SharedReg848_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg848_out;
SharedReg42_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg42_out;
   MUX_Product22_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg205_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg872_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg70_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg848_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg42_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_3_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_3_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product22_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_4_impl_out,
                 X => Delay1No258_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast);

SharedReg923_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg923_out;
SharedReg916_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg927_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg927_out;
SharedReg909_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product22_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg923_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_4_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_0_out,
                 Y => Delay1No258_out);

SharedReg809_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg809_out;
SharedReg61_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg241_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg241_out;
SharedReg95_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg95_out;
SharedReg874_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg874_out;
SharedReg72_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg72_out;
   MUX_Product22_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg809_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg241_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg95_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg874_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg72_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product22_4_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No260_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg75_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg924_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg924_out;
SharedReg64_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg64_out;
SharedReg209_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg76_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg76_out;
SharedReg932_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg932_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg924_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg64_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg76_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg932_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No260_out);

SharedReg909_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg739_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg739_out;
SharedReg916_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg866_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg866_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg739_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg866_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No262_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg932_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg932_out;
SharedReg77_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg924_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg924_out;
SharedReg67_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg67_out;
SharedReg199_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg199_out;
SharedReg67_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg67_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg932_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg924_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg67_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg199_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg67_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No262_out);

SharedReg868_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg868_out;
SharedReg909_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg743_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg743_out;
SharedReg916_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg868_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg743_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Product32_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_2_impl_out,
                 X => Delay1No264_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg69_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg932_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg932_out;
SharedReg79_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg79_out;
SharedReg924_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg924_out;
SharedReg56_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg56_out;
SharedReg202_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg202_out;
   MUX_Product32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg932_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg79_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg924_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg56_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg202_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_2_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_0_out,
                 Y => Delay1No264_out);

SharedReg913_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg870_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg870_out;
SharedReg909_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg804_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg804_out;
SharedReg916_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg870_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg804_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_2_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No266_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg221_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg82_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg932_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg932_out;
SharedReg81_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg81_out;
SharedReg924_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg924_out;
SharedReg58_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg58_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg932_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg81_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg924_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg58_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No266_out);

SharedReg912_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg872_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg872_out;
SharedReg909_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg805_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg805_out;
SharedReg916_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg872_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg805_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No268_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg924_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg924_out;
SharedReg73_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg73_out;
SharedReg257_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg257_out;
SharedReg97_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg97_out;
SharedReg932_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg932_out;
SharedReg83_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg83_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg924_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg73_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg257_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg97_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg932_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg83_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No268_out);

SharedReg755_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg755_out;
SharedReg916_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg874_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg874_out;
SharedReg909_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg755_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg874_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Subtract3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_0_impl_out,
                 X => Delay1No270_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg301_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg301_out;
SharedReg311_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg311_out;
SharedReg301_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg301_out;
SharedReg340_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg340_out;
SharedReg311_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg311_out;
SharedReg335_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg335_out;
   MUX_Subtract3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg301_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg311_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg301_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg340_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg311_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg335_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_0_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_0_out,
                 Y => Delay1No270_out);

Delay3No35_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast <= Delay3No35_out;
SharedReg345_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
SharedReg292_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg292_out;
SharedReg561_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg345_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg345_out;
SharedReg301_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg301_out;
   MUX_Subtract3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No35_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg292_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg345_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg301_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_0_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Subtract3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_1_impl_out,
                 X => Delay1No272_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg718_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg718_out;
SharedReg15_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg259_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg259_out;
SharedReg87_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg87_out;
SharedReg341_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg341_out;
SharedReg312_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg312_out;
   MUX_Subtract3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg718_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg259_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg87_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg341_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg312_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_1_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_0_out,
                 Y => Delay1No272_out);

Delay8No50_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast <= Delay8No50_out;
SharedReg31_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg87_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg87_out;
SharedReg541_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg541_out;
SharedReg563_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg563_out;
SharedReg346_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg346_out;
   MUX_Subtract3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay8No50_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg87_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg541_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg563_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg346_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_1_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Subtract3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_2_impl_out,
                 X => Delay1No274_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast);

SharedReg313_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg313_out;
SharedReg723_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg723_out;
SharedReg15_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg15_out;
SharedReg262_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg262_out;
SharedReg305_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg305_out;
SharedReg701_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg701_out;
   MUX_Subtract3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg313_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg723_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg15_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg262_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg305_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg701_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_2_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_2_impl_0_out,
                 Y => Delay1No274_out);

SharedReg347_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg347_out;
Delay8No51_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast <= Delay8No51_out;
SharedReg31_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg31_out;
SharedReg91_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg91_out;
SharedReg296_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg296_out;
SharedReg677_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg677_out;
   MUX_Subtract3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg347_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay8No51_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg31_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg91_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg296_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg677_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_2_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_2_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Subtract3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Subtract3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Subtract3_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_3_impl_out,
                 X => Delay1No276_out_to_Subtract3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Subtract3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg703_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg703_out;
SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg314_out;
SharedReg747_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg747_out;
SharedReg15_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg15_out;
SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg314_out;
SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg314_out;
   MUX_Subtract3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg703_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg747_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg15_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg314_out_to_MUX_Subtract3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_3_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_3_impl_0_out,
                 Y => Delay1No276_out);

SharedReg679_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg679_out;
SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg348_out;
Delay8No52_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_3_cast <= Delay8No52_out;
SharedReg31_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg31_out;
SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg348_out;
SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg348_out;
   MUX_Subtract3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg679_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay8No52_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg31_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg348_out_to_MUX_Subtract3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract3_3_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_3_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Product6_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_0_impl_out,
                 X => Delay1No278_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg919_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg919_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg925_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_0_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_0_out,
                 Y => Delay1No278_out);

SharedReg636_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg636_out;
SharedReg866_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg866_out;
SharedReg76_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg76_out;
SharedReg99_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg99_out;
SharedReg75_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg75_out;
SharedReg100_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg100_out;
   MUX_Product6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg636_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg866_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg76_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg99_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg75_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg100_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_0_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Product6_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_1_impl_out,
                 X => Delay1No280_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg919_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg925_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_1_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_0_out,
                 Y => Delay1No280_out);

SharedReg110_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg640_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg640_out;
SharedReg868_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg868_out;
SharedReg78_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg78_out;
SharedReg77_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg77_out;
SharedReg77_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg77_out;
   MUX_Product6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg640_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg868_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg78_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg77_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg77_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_1_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Product6_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_2_impl_out,
                 X => Delay1No282_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product6_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg919_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg925_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_2_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_2_impl_0_out,
                 Y => Delay1No282_out);

SharedReg79_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg112_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg726_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg726_out;
SharedReg870_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg870_out;
SharedReg69_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg69_out;
SharedReg79_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg79_out;
   MUX_Product6_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg726_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg870_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg69_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg79_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_2_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_2_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Product6_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_3_impl_out,
                 X => Delay1No284_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product6_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg919_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg925_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_3_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_0_out,
                 Y => Delay1No284_out);

SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg101_out;
SharedReg115_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg730_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg730_out;
SharedReg861_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg861_out;
SharedReg71_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg71_out;
   MUX_Product6_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg730_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg861_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg71_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_3_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Product6_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_4_impl_out,
                 X => Delay1No286_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg925_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg919_out;
   MUX_Product6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg925_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg919_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_4_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_0_out,
                 Y => Delay1No286_out);

SharedReg863_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg863_out;
SharedReg84_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg84_out;
SharedReg103_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg94_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg94_out;
SharedReg97_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg97_out;
SharedReg655_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg655_out;
   MUX_Product6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg863_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg84_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg94_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg97_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg655_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product6_4_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Product13_0_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Product13_0_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Product13_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_0_impl_out,
                 X => Delay1No288_out_to_Product13_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Product13_0_impl_parent_implementedSystem_port_1_cast);

SharedReg919_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product13_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg919_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg925_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product13_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_0_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_0_impl_0_out,
                 Y => Delay1No288_out);

SharedReg716_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg716_out;
SharedReg876_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg876_out;
SharedReg100_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg100_out;
SharedReg106_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg106_out;
SharedReg32_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg32_out;
SharedReg34_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg34_out;
   MUX_Product13_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg716_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg876_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg100_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg106_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg32_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg34_out_to_MUX_Product13_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_0_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_0_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Product13_1_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Product13_1_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Product13_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_1_impl_out,
                 X => Delay1No290_out_to_Product13_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Product13_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product13_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg919_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg925_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product13_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_1_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_1_impl_0_out,
                 Y => Delay1No290_out);

SharedReg89_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg721_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg721_out;
SharedReg878_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg878_out;
SharedReg110_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg110_out;
SharedReg109_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg109_out;
SharedReg35_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg35_out;
   MUX_Product13_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg721_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg878_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg109_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg35_out_to_MUX_Product13_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_1_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_1_impl_1_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Product13_2_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Product13_2_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Product13_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_2_impl_out,
                 X => Delay1No292_out_to_Product13_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Product13_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product13_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg919_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg925_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product13_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_2_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_2_impl_0_out,
                 Y => Delay1No292_out);

SharedReg38_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg151_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
SharedReg745_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg745_out;
SharedReg880_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg880_out;
SharedReg80_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg80_out;
SharedReg111_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg111_out;
   MUX_Product13_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg745_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg880_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg80_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg111_out_to_MUX_Product13_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_2_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_2_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Product13_3_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Product13_3_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Product13_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_3_impl_out,
                 X => Delay1No294_out_to_Product13_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Product13_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg919_out;
SharedReg925_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product13_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg919_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg925_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product13_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_3_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_3_impl_0_out,
                 Y => Delay1No294_out);

SharedReg114_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg57_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg57_out;
SharedReg156_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg156_out;
SharedReg749_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg749_out;
SharedReg872_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg872_out;
SharedReg82_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg82_out;
   MUX_Product13_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg57_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg156_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg749_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg872_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg82_out_to_MUX_Product13_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_3_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_3_impl_1_out,
                 Y => Delay1No295_out);

Delay1No296_out_to_Product13_4_impl_parent_implementedSystem_port_0_cast <= Delay1No296_out;
Delay1No297_out_to_Product13_4_impl_parent_implementedSystem_port_1_cast <= Delay1No297_out;
   Product13_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_4_impl_out,
                 X => Delay1No296_out_to_Product13_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No297_out_to_Product13_4_impl_parent_implementedSystem_port_1_cast);

SharedReg925_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg925_out;
SharedReg906_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg902_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg919_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg919_out;
   MUX_Product13_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg925_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg919_out_to_MUX_Product13_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_4_impl_0_out);

   Delay1No296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_4_impl_0_out,
                 Y => Delay1No296_out);

SharedReg874_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg874_out;
SharedReg95_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg116_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg60_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg62_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg62_out;
SharedReg734_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg734_out;
   MUX_Product13_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg874_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg116_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg62_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg734_out_to_MUX_Product13_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product13_4_impl_1_out);

   Delay1No297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_4_impl_1_out,
                 Y => Delay1No297_out);

Delay1No298_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No298_out;
Delay1No299_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No299_out;
   Product23_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_0_impl_out,
                 X => Delay1No298_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No299_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg921_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg921_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg930_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_0_impl_0_out);

   Delay1No298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_0_out,
                 Y => Delay1No298_out);

SharedReg636_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg636_out;
SharedReg866_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg866_out;
SharedReg76_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg76_out;
SharedReg99_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg99_out;
SharedReg75_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg75_out;
SharedReg100_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg100_out;
   MUX_Product23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg636_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg866_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg76_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg99_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg75_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg100_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_0_impl_1_out);

   Delay1No299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_1_out,
                 Y => Delay1No299_out);

Delay1No300_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No300_out;
Delay1No301_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No301_out;
   Product23_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_1_impl_out,
                 X => Delay1No300_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No301_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg918_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg921_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg930_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_1_impl_0_out);

   Delay1No300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_0_out,
                 Y => Delay1No300_out);

SharedReg110_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg640_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg640_out;
SharedReg868_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg868_out;
SharedReg78_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg78_out;
SharedReg77_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg77_out;
SharedReg77_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg77_out;
   MUX_Product23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg640_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg868_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg78_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg77_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg77_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_1_impl_1_out);

   Delay1No301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_1_out,
                 Y => Delay1No301_out);

Delay1No302_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No302_out;
Delay1No303_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No303_out;
   Product23_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_2_impl_out,
                 X => Delay1No302_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No303_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg921_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg930_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_2_impl_0_out);

   Delay1No302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_0_out,
                 Y => Delay1No302_out);

SharedReg79_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg79_out;
SharedReg112_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg726_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg726_out;
SharedReg870_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg870_out;
SharedReg69_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg69_out;
SharedReg79_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg79_out;
   MUX_Product23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg79_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg726_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg870_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg69_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg79_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_2_impl_1_out);

   Delay1No303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_1_out,
                 Y => Delay1No303_out);

Delay1No304_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast <= Delay1No304_out;
Delay1No305_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast <= Delay1No305_out;
   Product23_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_3_impl_out,
                 X => Delay1No304_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No305_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast);

SharedReg912_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product23_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg921_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg930_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_3_impl_0_out);

   Delay1No304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_0_out,
                 Y => Delay1No304_out);

SharedReg101_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg101_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg101_out;
SharedReg115_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg730_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg730_out;
SharedReg861_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg861_out;
SharedReg71_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg71_out;
   MUX_Product23_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg730_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg861_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg71_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_3_impl_1_out);

   Delay1No305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_1_out,
                 Y => Delay1No305_out);

Delay1No306_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast <= Delay1No306_out;
Delay1No307_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast <= Delay1No307_out;
   Product23_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_4_impl_out,
                 X => Delay1No306_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No307_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast);

SharedReg930_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg921_out;
   MUX_Product23_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg930_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg921_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_4_impl_0_out);

   Delay1No306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_0_out,
                 Y => Delay1No306_out);

SharedReg863_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg863_out;
SharedReg84_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg84_out;
SharedReg103_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg94_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg94_out;
SharedReg97_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg97_out;
SharedReg655_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg655_out;
   MUX_Product23_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg863_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg84_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg94_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg97_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg655_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product23_4_impl_1_out);

   Delay1No307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_1_out,
                 Y => Delay1No307_out);

Delay1No308_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No308_out;
Delay1No309_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No309_out;
   Product33_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_0_impl_out,
                 X => Delay1No308_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No309_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg716_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg716_out;
SharedReg876_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg876_out;
SharedReg100_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg100_out;
SharedReg106_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg106_out;
SharedReg32_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg32_out;
SharedReg34_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg34_out;
   MUX_Product33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg716_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg876_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg100_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg106_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg32_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg34_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_0_impl_0_out);

   Delay1No308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_0_out,
                 Y => Delay1No308_out);

SharedReg921_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg921_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg930_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_0_impl_1_out);

   Delay1No309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_1_out,
                 Y => Delay1No309_out);

Delay1No310_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast <= Delay1No310_out;
Delay1No311_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast <= Delay1No311_out;
   Product33_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_1_impl_out,
                 X => Delay1No310_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No311_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg721_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg721_out;
SharedReg878_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg878_out;
SharedReg110_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg110_out;
SharedReg109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg109_out;
SharedReg35_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg35_out;
   MUX_Product33_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg721_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg878_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg109_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg35_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_1_impl_0_out);

   Delay1No310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_0_out,
                 Y => Delay1No310_out);

SharedReg918_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product33_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg921_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg930_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_1_impl_1_out);

   Delay1No311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_1_out,
                 Y => Delay1No311_out);

Delay1No312_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast <= Delay1No312_out;
Delay1No313_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast <= Delay1No313_out;
   Product33_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_2_impl_out,
                 X => Delay1No312_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No313_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast);

SharedReg38_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg151_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg151_out;
SharedReg745_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg745_out;
SharedReg880_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg880_out;
SharedReg80_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg80_out;
SharedReg111_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg111_out;
   MUX_Product33_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg745_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg880_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg80_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg111_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_2_impl_0_out);

   Delay1No312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_0_out,
                 Y => Delay1No312_out);

SharedReg913_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product33_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg921_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg930_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_2_impl_1_out);

   Delay1No313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_1_out,
                 Y => Delay1No313_out);

Delay1No314_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast <= Delay1No314_out;
Delay1No315_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast <= Delay1No315_out;
   Product33_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_3_impl_out,
                 X => Delay1No314_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No315_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast);

SharedReg114_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg57_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg57_out;
SharedReg156_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg156_out;
SharedReg749_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg749_out;
SharedReg872_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg872_out;
SharedReg82_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg82_out;
   MUX_Product33_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg57_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg156_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg749_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg872_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg82_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_3_impl_0_out);

   Delay1No314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_0_out,
                 Y => Delay1No314_out);

SharedReg912_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg921_out;
SharedReg930_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product33_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg921_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg930_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_3_impl_1_out);

   Delay1No315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_1_out,
                 Y => Delay1No315_out);

Delay1No316_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast <= Delay1No316_out;
Delay1No317_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast <= Delay1No317_out;
   Product33_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_4_impl_out,
                 X => Delay1No316_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No317_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast);

SharedReg874_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg874_out;
SharedReg95_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg116_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg60_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
SharedReg62_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg62_out;
SharedReg734_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg734_out;
   MUX_Product33_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg874_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg116_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg62_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg734_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_4_impl_0_out);

   Delay1No316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_0_out,
                 Y => Delay1No316_out);

SharedReg930_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg930_out;
SharedReg916_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg912_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg921_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg921_out;
   MUX_Product33_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg930_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg921_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product33_4_impl_1_out);

   Delay1No317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_1_out,
                 Y => Delay1No317_out);

Delay1No318_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No318_out;
Delay1No319_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No319_out;
   Subtract4_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_1_impl_out,
                 X => Delay1No318_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No319_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg336_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg336_out;
SharedReg303_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg303_out;
SharedReg312_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg312_out;
SharedReg303_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg303_out;
SharedReg699_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg699_out;
SharedReg364_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg364_out;
   MUX_Subtract4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg336_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg303_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg312_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg303_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg699_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg364_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_1_impl_0_out);

   Delay1No318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_0_out,
                 Y => Delay1No318_out);

SharedReg303_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg303_out;
Delay3No36_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast <= Delay3No36_out;
SharedReg346_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg294_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg294_out;
SharedReg675_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg675_out;
SharedReg379_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg379_out;
   MUX_Subtract4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg303_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No36_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg346_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg675_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg379_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_1_impl_1_out);

   Delay1No319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_1_out,
                 Y => Delay1No319_out);

Delay1No320_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No320_out;
Delay1No321_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No321_out;
   Subtract4_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_2_impl_out,
                 X => Delay1No320_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No321_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg365_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg365_out;
SharedReg337_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg337_out;
SharedReg305_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg305_out;
SharedReg313_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg313_out;
SharedReg313_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg313_out;
SharedReg763_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg763_out;
   MUX_Subtract4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg365_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg337_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg305_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg313_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg313_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg763_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_2_impl_0_out);

   Delay1No320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_0_out,
                 Y => Delay1No320_out);

SharedReg380_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg380_out;
SharedReg305_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg305_out;
Delay3No37_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast <= Delay3No37_out;
SharedReg347_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg347_out;
SharedReg347_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg347_out;
SharedReg772_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg772_out;
   MUX_Subtract4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg380_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg305_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No37_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg347_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg347_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg772_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_2_impl_1_out);

   Delay1No321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_1_out,
                 Y => Delay1No321_out);

Delay1No322_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No322_out;
Delay1No323_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No323_out;
   Subtract4_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_3_impl_out,
                 X => Delay1No322_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No323_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg765_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg765_out;
SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg366_out;
SharedReg338_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg307_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg307_out;
SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg366_out;
SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg366_out;
   MUX_Subtract4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg765_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg338_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg307_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg366_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_3_impl_0_out);

   Delay1No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_0_out,
                 Y => Delay1No322_out);

SharedReg774_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg774_out;
SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg381_out;
SharedReg307_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg307_out;
Delay3No38_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast <= Delay3No38_out;
SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg381_out;
SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg381_out;
   MUX_Subtract4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg774_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg307_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No38_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg381_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_3_impl_1_out);

   Delay1No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_1_out,
                 Y => Delay1No323_out);

Delay1No324_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No324_out;
Delay1No325_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No325_out;
   Subtract4_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_4_impl_out,
                 X => Delay1No324_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No325_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg423_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg423_out;
SharedReg767_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg767_out;
SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg367_out;
SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg367_out;
SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg367_out;
   MUX_Subtract4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg423_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg767_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg367_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_4_impl_0_out);

   Delay1No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_0_out,
                 Y => Delay1No324_out);

SharedReg16_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg472_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg472_out;
SharedReg776_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg776_out;
SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg382_out;
SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg382_out;
SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg382_out;
   MUX_Subtract4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg472_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg776_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg382_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract4_4_impl_1_out);

   Delay1No325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_1_out,
                 Y => Delay1No325_out);

Delay1No326_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast <= Delay1No326_out;
Delay1No327_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast <= Delay1No327_out;
   Subtract5_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract5_4_impl_out,
                 X => Delay1No326_out_to_Subtract5_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No327_out_to_Subtract5_4_impl_parent_implementedSystem_port_1_cast);

SharedReg367_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg315_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg315_out;
SharedReg344_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg344_out;
SharedReg806_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg806_out;
SharedReg339_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg339_out;
SharedReg315_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg315_out;
   MUX_Subtract5_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg315_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg344_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg806_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg339_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg315_out_to_MUX_Subtract5_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract5_4_impl_0_out);

   Delay1No326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_4_impl_0_out,
                 Y => Delay1No326_out);

SharedReg382_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg382_out;
SharedReg349_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg349_out;
SharedReg569_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg569_out;
Delay8No53_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast <= Delay8No53_out;
SharedReg309_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg309_out;
SharedReg349_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg349_out;
   MUX_Subtract5_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg382_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg349_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg569_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay8No53_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg309_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg349_out_to_MUX_Subtract5_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract5_4_impl_1_out);

   Delay1No327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_4_impl_1_out,
                 Y => Delay1No327_out);

Delay1No328_out_to_Subtract6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No328_out;
Delay1No329_out_to_Subtract6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No329_out;
   Subtract6_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_0_impl_out,
                 X => Delay1No328_out_to_Subtract6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No329_out_to_Subtract6_0_impl_parent_implementedSystem_port_1_cast);

Delay4No50_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No50_out;
SharedReg663_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg663_out;
SharedReg363_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg363_out;
SharedReg759_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg759_out;
SharedReg480_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg480_out;
SharedReg363_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg363_out;
   MUX_Subtract6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No50_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg663_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg363_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg759_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg480_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg363_out_to_MUX_Subtract6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_0_impl_0_out);

   Delay1No328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_0_impl_0_out,
                 Y => Delay1No328_out);

Delay4No65_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No65_out;
SharedReg688_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg688_out;
SharedReg378_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg378_out;
SharedReg768_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg768_out;
SharedReg510_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg510_out;
SharedReg378_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg378_out;
   MUX_Subtract6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No65_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg688_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg378_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg768_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg510_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg378_out_to_MUX_Subtract6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_0_impl_1_out);

   Delay1No329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_0_impl_1_out,
                 Y => Delay1No329_out);

Delay1No330_out_to_Subtract6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No330_out;
Delay1No331_out_to_Subtract6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No331_out;
   Subtract6_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_1_impl_out,
                 X => Delay1No330_out_to_Subtract6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No331_out_to_Subtract6_1_impl_parent_implementedSystem_port_1_cast);

SharedReg364_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg364_out;
Delay4No51_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No51_out;
SharedReg665_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg665_out;
SharedReg364_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg364_out;
SharedReg416_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg416_out;
SharedReg552_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg552_out;
   MUX_Subtract6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg364_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No51_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg665_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg364_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg416_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg552_out_to_MUX_Subtract6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_1_impl_0_out);

   Delay1No330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_1_impl_0_out,
                 Y => Delay1No330_out);

SharedReg379_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg379_out;
Delay4No66_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No66_out;
SharedReg689_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg689_out;
SharedReg379_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg465_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg465_out;
SharedReg587_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg587_out;
   MUX_Subtract6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No66_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg689_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg465_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg587_out_to_MUX_Subtract6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_1_impl_1_out);

   Delay1No331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_1_impl_1_out,
                 Y => Delay1No331_out);

Delay1No332_out_to_Subtract6_2_impl_parent_implementedSystem_port_0_cast <= Delay1No332_out;
Delay1No333_out_to_Subtract6_2_impl_parent_implementedSystem_port_1_cast <= Delay1No333_out;
   Subtract6_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_2_impl_out,
                 X => Delay1No332_out_to_Subtract6_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No333_out_to_Subtract6_2_impl_parent_implementedSystem_port_1_cast);

SharedReg554_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg554_out;
SharedReg365_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg365_out;
Delay4No52_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_3_cast <= Delay4No52_out;
SharedReg667_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg667_out;
SharedReg419_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg419_out;
SharedReg782_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg782_out;
   MUX_Subtract6_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg554_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg365_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No52_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg667_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg419_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg782_out_to_MUX_Subtract6_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_2_impl_0_out);

   Delay1No332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_2_impl_0_out,
                 Y => Delay1No332_out);

SharedReg589_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg589_out;
SharedReg380_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg380_out;
Delay4No67_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No67_out;
SharedReg690_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg690_out;
SharedReg468_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg468_out;
SharedReg793_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg793_out;
   MUX_Subtract6_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg589_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg380_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No67_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg690_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg468_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg793_out_to_MUX_Subtract6_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_2_impl_1_out);

   Delay1No333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_2_impl_1_out,
                 Y => Delay1No333_out);

Delay1No334_out_to_Subtract6_3_impl_parent_implementedSystem_port_0_cast <= Delay1No334_out;
Delay1No335_out_to_Subtract6_3_impl_parent_implementedSystem_port_1_cast <= Delay1No335_out;
   Subtract6_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract6_3_impl_out,
                 X => Delay1No334_out_to_Subtract6_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No335_out_to_Subtract6_3_impl_parent_implementedSystem_port_1_cast);

SharedReg784_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg784_out;
SharedReg556_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg366_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg366_out;
Delay4No53_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_4_cast <= Delay4No53_out;
SharedReg_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg420_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg420_out;
   MUX_Subtract6_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg784_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg366_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No53_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg420_out_to_MUX_Subtract6_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_3_impl_0_out);

   Delay1No334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_3_impl_0_out,
                 Y => Delay1No334_out);

SharedReg795_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg795_out;
SharedReg591_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg591_out;
SharedReg381_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg381_out;
Delay4No68_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_4_cast <= Delay4No68_out;
SharedReg16_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg469_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg469_out;
   MUX_Subtract6_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg795_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg591_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg381_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No68_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg469_out_to_MUX_Subtract6_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract6_3_impl_1_out);

   Delay1No335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract6_3_impl_1_out,
                 Y => Delay1No335_out);

Delay1No336_out_to_Product9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No336_out;
Delay1No337_out_to_Product9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No337_out;
   Product9_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_0_impl_out,
                 X => Delay1No336_out_to_Product9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No337_out_to_Product9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg935_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg935_out;
SharedReg936_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg936_out;
SharedReg929_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg935_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg936_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_0_impl_0_out);

   Delay1No336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_0_impl_0_out,
                 Y => Delay1No336_out);

SharedReg885_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg885_out;
SharedReg812_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg812_out;
SharedReg886_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg886_out;
SharedReg119_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg119_out;
SharedReg717_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg717_out;
SharedReg65_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg65_out;
   MUX_Product9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg885_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg812_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg886_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg119_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg717_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg65_out_to_MUX_Product9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_0_impl_1_out);

   Delay1No337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_0_impl_1_out,
                 Y => Delay1No337_out);

Delay1No338_out_to_Product9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No338_out;
Delay1No339_out_to_Product9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No339_out;
   Product9_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_1_impl_out,
                 X => Delay1No338_out_to_Product9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No339_out_to_Product9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg935_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg935_out;
SharedReg936_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg936_out;
SharedReg929_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg935_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg936_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_1_impl_0_out);

   Delay1No338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_1_impl_0_out,
                 Y => Delay1No338_out);

SharedReg54_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg887_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg887_out;
SharedReg815_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg815_out;
SharedReg888_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg888_out;
SharedReg122_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg122_out;
SharedReg641_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg641_out;
   MUX_Product9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg887_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg815_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg888_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg122_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg641_out_to_MUX_Product9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_1_impl_1_out);

   Delay1No339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_1_impl_1_out,
                 Y => Delay1No339_out);

Delay1No340_out_to_Product9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No340_out;
Delay1No341_out_to_Product9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No341_out;
   Product9_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_2_impl_out,
                 X => Delay1No340_out_to_Product9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No341_out_to_Product9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg935_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg935_out;
SharedReg936_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg936_out;
SharedReg929_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg935_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg936_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product9_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_2_impl_0_out);

   Delay1No340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_2_impl_0_out,
                 Y => Delay1No340_out);

SharedReg727_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg727_out;
SharedReg40_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg889_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg889_out;
SharedReg818_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg818_out;
SharedReg880_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg880_out;
SharedReg125_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg125_out;
   MUX_Product9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg727_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg889_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg818_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg880_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg125_out_to_MUX_Product9_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_2_impl_1_out);

   Delay1No341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_2_impl_1_out,
                 Y => Delay1No341_out);

Delay1No342_out_to_Product9_3_impl_parent_implementedSystem_port_0_cast <= Delay1No342_out;
Delay1No343_out_to_Product9_3_impl_parent_implementedSystem_port_1_cast <= Delay1No343_out;
   Product9_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_3_impl_out,
                 X => Delay1No342_out_to_Product9_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No343_out_to_Product9_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg935_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg935_out;
SharedReg936_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg936_out;
SharedReg929_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product9_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg935_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg936_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product9_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_3_impl_0_out);

   Delay1No342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_3_impl_0_out,
                 Y => Delay1No342_out);

SharedReg127_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg750_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg750_out;
SharedReg59_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg881_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg881_out;
SharedReg892_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg892_out;
SharedReg872_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg872_out;
   MUX_Product9_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg750_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg59_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg881_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg892_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg872_out_to_MUX_Product9_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_3_impl_1_out);

   Delay1No343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_3_impl_1_out,
                 Y => Delay1No343_out);

Delay1No344_out_to_Product9_4_impl_parent_implementedSystem_port_0_cast <= Delay1No344_out;
Delay1No345_out_to_Product9_4_impl_parent_implementedSystem_port_1_cast <= Delay1No345_out;
   Product9_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product9_4_impl_out,
                 X => Delay1No344_out_to_Product9_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No345_out_to_Product9_4_impl_parent_implementedSystem_port_1_cast);

SharedReg936_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg936_out;
SharedReg929_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg935_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg935_out;
   MUX_Product9_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg936_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg935_out_to_MUX_Product9_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_4_impl_0_out);

   Delay1No344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_4_impl_0_out,
                 Y => Delay1No344_out);

SharedReg825_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg825_out;
SharedReg884_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg884_out;
SharedReg130_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg130_out;
SharedReg809_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg809_out;
SharedReg85_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg85_out;
SharedReg883_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg883_out;
   MUX_Product9_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg825_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg884_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg130_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg809_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg85_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg883_out_to_MUX_Product9_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product9_4_impl_1_out);

   Delay1No345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product9_4_impl_1_out,
                 Y => Delay1No345_out);

Delay1No346_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast <= Delay1No346_out;
Delay1No347_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast <= Delay1No347_out;
   Product26_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_0_impl_out,
                 X => Delay1No346_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No347_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast);

SharedReg937_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg937_out;
SharedReg812_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg812_out;
SharedReg929_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product26_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg937_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg812_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_0_impl_0_out);

   Delay1No346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_0_out,
                 Y => Delay1No346_out);

SharedReg885_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg885_out;
SharedReg938_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg938_out;
SharedReg812_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg812_out;
SharedReg133_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg133_out;
SharedReg739_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg739_out;
SharedReg163_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg163_out;
   MUX_Product26_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg885_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg938_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg812_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg133_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg163_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_0_impl_1_out);

   Delay1No347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_1_out,
                 Y => Delay1No347_out);

Delay1No348_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No348_out;
Delay1No349_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No349_out;
   Product26_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_1_impl_out,
                 X => Delay1No348_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No349_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg937_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg937_out;
SharedReg815_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg815_out;
SharedReg929_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg937_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg815_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_1_impl_0_out);

   Delay1No348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_0_out,
                 Y => Delay1No348_out);

SharedReg166_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg887_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg887_out;
SharedReg938_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg938_out;
SharedReg815_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg815_out;
SharedReg136_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg136_out;
SharedReg722_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg722_out;
   MUX_Product26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg887_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg938_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg815_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg136_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg722_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_1_impl_1_out);

   Delay1No349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_1_out,
                 Y => Delay1No349_out);

Delay1No350_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast <= Delay1No350_out;
Delay1No351_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast <= Delay1No351_out;
   Product26_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_2_impl_out,
                 X => Delay1No350_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No351_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg937_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg937_out;
SharedReg818_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg818_out;
SharedReg929_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product26_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg937_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg818_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_2_impl_0_out);

   Delay1No350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_2_impl_0_out,
                 Y => Delay1No350_out);

SharedReg746_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg746_out;
SharedReg169_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg169_out;
SharedReg889_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg889_out;
SharedReg938_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg938_out;
SharedReg890_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg890_out;
SharedReg139_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg139_out;
   MUX_Product26_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg746_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg169_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg889_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg938_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg890_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_2_impl_1_out);

   Delay1No351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_2_impl_1_out,
                 Y => Delay1No351_out);

Delay1No352_out_to_Product26_3_impl_parent_implementedSystem_port_0_cast <= Delay1No352_out;
Delay1No353_out_to_Product26_3_impl_parent_implementedSystem_port_1_cast <= Delay1No353_out;
   Product26_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_3_impl_out,
                 X => Delay1No352_out_to_Product26_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No353_out_to_Product26_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg937_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg937_out;
SharedReg892_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg892_out;
SharedReg929_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product26_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg937_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg892_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product26_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_3_impl_0_out);

   Delay1No352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_3_impl_0_out,
                 Y => Delay1No352_out);

SharedReg142_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg805_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg805_out;
SharedReg144_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg144_out;
SharedReg881_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg881_out;
SharedReg938_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg938_out;
SharedReg882_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg882_out;
   MUX_Product26_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg805_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg144_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg881_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg938_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg882_out_to_MUX_Product26_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_3_impl_1_out);

   Delay1No353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_3_impl_1_out,
                 Y => Delay1No353_out);

Delay1No354_out_to_Product26_4_impl_parent_implementedSystem_port_0_cast <= Delay1No354_out;
Delay1No355_out_to_Product26_4_impl_parent_implementedSystem_port_1_cast <= Delay1No355_out;
   Product26_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_4_impl_out,
                 X => Delay1No354_out_to_Product26_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No355_out_to_Product26_4_impl_parent_implementedSystem_port_1_cast);

SharedReg825_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg825_out;
SharedReg929_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg903_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg937_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg937_out;
   MUX_Product26_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg825_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg937_out_to_MUX_Product26_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_4_impl_0_out);

   Delay1No354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_4_impl_0_out,
                 Y => Delay1No354_out);

SharedReg938_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg938_out;
SharedReg825_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg825_out;
SharedReg145_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg145_out;
SharedReg863_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg863_out;
SharedReg132_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg132_out;
SharedReg883_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg883_out;
   MUX_Product26_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg938_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg825_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg145_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg863_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg132_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg883_out_to_MUX_Product26_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product26_4_impl_1_out);

   Delay1No355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_4_impl_1_out,
                 Y => Delay1No355_out);

Delay1No356_out_to_Subtract7_0_impl_parent_implementedSystem_port_0_cast <= Delay1No356_out;
Delay1No357_out_to_Subtract7_0_impl_parent_implementedSystem_port_1_cast <= Delay1No357_out;
   Subtract7_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_0_impl_out,
                 X => Delay1No356_out_to_Subtract7_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No357_out_to_Subtract7_0_impl_parent_implementedSystem_port_1_cast);

SharedReg363_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg363_out;
SharedReg_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg415_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg414_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg414_out;
SharedReg550_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg550_out;
SharedReg415_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg415_out;
   MUX_Subtract7_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg363_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg415_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg414_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg550_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg415_out_to_MUX_Subtract7_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_0_impl_0_out);

   Delay1No356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_0_impl_0_out,
                 Y => Delay1No356_out);

SharedReg378_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg378_out;
SharedReg16_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg464_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg464_out;
SharedReg463_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg463_out;
SharedReg585_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg585_out;
SharedReg424_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg424_out;
   MUX_Subtract7_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg378_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg464_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg463_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg585_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg424_out_to_MUX_Subtract7_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_0_impl_1_out);

   Delay1No357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_0_impl_1_out,
                 Y => Delay1No357_out);

Delay1No358_out_to_Subtract7_1_impl_parent_implementedSystem_port_0_cast <= Delay1No358_out;
Delay1No359_out_to_Subtract7_1_impl_parent_implementedSystem_port_1_cast <= Delay1No359_out;
   Subtract7_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_1_impl_out,
                 X => Delay1No358_out_to_Subtract7_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No359_out_to_Subtract7_1_impl_parent_implementedSystem_port_1_cast);

SharedReg417_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg417_out;
SharedReg364_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg364_out;
SharedReg_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg_out;
SharedReg417_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg417_out;
SharedReg780_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg780_out;
SharedReg684_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg684_out;
   MUX_Subtract7_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg417_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg364_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg417_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg780_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg684_out_to_MUX_Subtract7_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_1_impl_0_out);

   Delay1No358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_1_impl_0_out,
                 Y => Delay1No358_out);

SharedReg426_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg426_out;
SharedReg379_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg379_out;
SharedReg16_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg466_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg466_out;
SharedReg791_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg791_out;
SharedReg708_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg708_out;
   MUX_Subtract7_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg426_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg379_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg466_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg791_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg708_out_to_MUX_Subtract7_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_1_impl_1_out);

   Delay1No359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_1_impl_1_out,
                 Y => Delay1No359_out);

Delay1No360_out_to_Subtract7_2_impl_parent_implementedSystem_port_0_cast <= Delay1No360_out;
Delay1No361_out_to_Subtract7_2_impl_parent_implementedSystem_port_1_cast <= Delay1No361_out;
   Subtract7_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_2_impl_out,
                 X => Delay1No360_out_to_Subtract7_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No361_out_to_Subtract7_2_impl_parent_implementedSystem_port_1_cast);

SharedReg685_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg685_out;
SharedReg419_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg419_out;
SharedReg365_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg365_out;
SharedReg_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg_out;
SharedReg418_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg418_out;
SharedReg197_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg197_out;
   MUX_Subtract7_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg685_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg419_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg365_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg418_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Subtract7_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_2_impl_0_out);

   Delay1No360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_2_impl_0_out,
                 Y => Delay1No360_out);

SharedReg710_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg710_out;
SharedReg428_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg428_out;
SharedReg380_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg380_out;
SharedReg16_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg16_out;
SharedReg467_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg467_out;
SharedReg203_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg203_out;
   MUX_Subtract7_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg710_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg428_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg380_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg16_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg467_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg203_out_to_MUX_Subtract7_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_2_impl_1_out);

   Delay1No361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_2_impl_1_out,
                 Y => Delay1No361_out);

Delay1No362_out_to_Subtract7_3_impl_parent_implementedSystem_port_0_cast <= Delay1No362_out;
Delay1No363_out_to_Subtract7_3_impl_parent_implementedSystem_port_1_cast <= Delay1No363_out;
   Subtract7_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_3_impl_out,
                 X => Delay1No362_out_to_Subtract7_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No363_out_to_Subtract7_3_impl_parent_implementedSystem_port_1_cast);

SharedReg184_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg686_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg686_out;
SharedReg421_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg421_out;
SharedReg366_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg366_out;
SharedReg1_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg487_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg487_out;
   MUX_Subtract7_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg686_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg421_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg366_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg487_out_to_MUX_Subtract7_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_3_impl_0_out);

   Delay1No362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_3_impl_0_out,
                 Y => Delay1No362_out);

SharedReg222_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg222_out;
SharedReg712_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg712_out;
SharedReg430_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg430_out;
SharedReg381_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg381_out;
SharedReg17_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg17_out;
SharedReg517_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg517_out;
   MUX_Subtract7_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg222_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg712_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg430_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg381_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg17_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg517_out_to_MUX_Subtract7_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_3_impl_1_out);

   Delay1No363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_3_impl_1_out,
                 Y => Delay1No363_out);

Delay1No364_out_to_Subtract7_4_impl_parent_implementedSystem_port_0_cast <= Delay1No364_out;
Delay1No365_out_to_Subtract7_4_impl_parent_implementedSystem_port_1_cast <= Delay1No365_out;
   Subtract7_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract7_4_impl_out,
                 X => Delay1No364_out_to_Subtract7_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No365_out_to_Subtract7_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg422_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg422_out;
SharedReg488_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg488_out;
SharedReg423_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg423_out;
Delay4No74_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_6_cast <= Delay4No74_out;
   MUX_Subtract7_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg422_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg422_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg488_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No74_out_to_MUX_Subtract7_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_4_impl_0_out);

   Delay1No364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_4_impl_0_out,
                 Y => Delay1No364_out);

SharedReg17_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg17_out;
SharedReg471_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg471_out;
SharedReg471_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg471_out;
SharedReg518_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg518_out;
SharedReg432_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg432_out;
Delay4No89_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_6_cast <= Delay4No89_out;
   MUX_Subtract7_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg17_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg471_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg471_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg518_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg432_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay4No89_out_to_MUX_Subtract7_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract7_4_impl_1_out);

   Delay1No365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract7_4_impl_1_out,
                 Y => Delay1No365_out);

Delay1No366_out_to_Product17_0_impl_parent_implementedSystem_port_0_cast <= Delay1No366_out;
Delay1No367_out_to_Product17_0_impl_parent_implementedSystem_port_1_cast <= Delay1No367_out;
   Product17_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_0_impl_out,
                 X => Delay1No366_out_to_Product17_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No367_out_to_Product17_0_impl_parent_implementedSystem_port_1_cast);

SharedReg939_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg939_out;
SharedReg900_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product17_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg939_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product17_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_0_impl_0_out);

   Delay1No366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_0_impl_0_out,
                 Y => Delay1No366_out);

SharedReg849_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg134_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg134_out;
SharedReg886_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg886_out;
SharedReg119_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg119_out;
SharedReg717_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg717_out;
SharedReg65_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg65_out;
   MUX_Product17_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg886_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg119_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg717_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg65_out_to_MUX_Product17_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_0_impl_1_out);

   Delay1No367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_0_impl_1_out,
                 Y => Delay1No367_out);

Delay1No368_out_to_Product17_1_impl_parent_implementedSystem_port_0_cast <= Delay1No368_out;
Delay1No369_out_to_Product17_1_impl_parent_implementedSystem_port_1_cast <= Delay1No369_out;
   Product17_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_1_impl_out,
                 X => Delay1No368_out_to_Product17_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No369_out_to_Product17_1_impl_parent_implementedSystem_port_1_cast);

SharedReg918_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg939_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg939_out;
SharedReg900_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product17_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg939_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product17_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_1_impl_0_out);

   Delay1No368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_1_impl_0_out,
                 Y => Delay1No368_out);

SharedReg54_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg851_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg851_out;
SharedReg159_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg159_out;
SharedReg888_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg888_out;
SharedReg122_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg122_out;
SharedReg641_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg641_out;
   MUX_Product17_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg851_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg159_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg888_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg122_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg641_out_to_MUX_Product17_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_1_impl_1_out);

   Delay1No369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_1_impl_1_out,
                 Y => Delay1No369_out);

Delay1No370_out_to_Product17_2_impl_parent_implementedSystem_port_0_cast <= Delay1No370_out;
Delay1No371_out_to_Product17_2_impl_parent_implementedSystem_port_1_cast <= Delay1No371_out;
   Product17_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_2_impl_out,
                 X => Delay1No370_out_to_Product17_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No371_out_to_Product17_2_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg939_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg939_out;
SharedReg900_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product17_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg939_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product17_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_2_impl_0_out);

   Delay1No370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_2_impl_0_out,
                 Y => Delay1No370_out);

SharedReg727_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg727_out;
SharedReg40_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg853_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg853_out;
SharedReg168_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
SharedReg880_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg880_out;
SharedReg125_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg125_out;
   MUX_Product17_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg727_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg853_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg880_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg125_out_to_MUX_Product17_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_2_impl_1_out);

   Delay1No371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_2_impl_1_out,
                 Y => Delay1No371_out);

Delay1No372_out_to_Product17_3_impl_parent_implementedSystem_port_0_cast <= Delay1No372_out;
Delay1No373_out_to_Product17_3_impl_parent_implementedSystem_port_1_cast <= Delay1No373_out;
   Product17_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_3_impl_out,
                 X => Delay1No372_out_to_Product17_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No373_out_to_Product17_3_impl_parent_implementedSystem_port_1_cast);

SharedReg912_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg939_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg939_out;
SharedReg900_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product17_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg939_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product17_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_3_impl_0_out);

   Delay1No372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_3_impl_0_out,
                 Y => Delay1No372_out);

SharedReg127_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg750_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg750_out;
SharedReg59_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg840_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg840_out;
SharedReg143_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg143_out;
SharedReg872_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg872_out;
   MUX_Product17_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg750_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg59_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg840_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg143_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg872_out_to_MUX_Product17_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_3_impl_1_out);

   Delay1No373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_3_impl_1_out,
                 Y => Delay1No373_out);

Delay1No374_out_to_Product17_4_impl_parent_implementedSystem_port_0_cast <= Delay1No374_out;
Delay1No375_out_to_Product17_4_impl_parent_implementedSystem_port_1_cast <= Delay1No375_out;
   Product17_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_4_impl_out,
                 X => Delay1No374_out_to_Product17_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No375_out_to_Product17_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg939_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg939_out;
   MUX_Product17_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg939_out_to_MUX_Product17_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_4_impl_0_out);

   Delay1No374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_4_impl_0_out,
                 Y => Delay1No374_out);

SharedReg117_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg884_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg884_out;
SharedReg130_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg130_out;
SharedReg809_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg809_out;
SharedReg85_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg85_out;
SharedReg856_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg856_out;
   MUX_Product17_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg884_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg130_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg809_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg85_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg856_out_to_MUX_Product17_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product17_4_impl_1_out);

   Delay1No375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_4_impl_1_out,
                 Y => Delay1No375_out);

Delay1No376_out_to_Product37_0_impl_parent_implementedSystem_port_0_cast <= Delay1No376_out;
Delay1No377_out_to_Product37_0_impl_parent_implementedSystem_port_1_cast <= Delay1No377_out;
   Product37_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_0_impl_out,
                 X => Delay1No376_out_to_Product37_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No377_out_to_Product37_0_impl_parent_implementedSystem_port_1_cast);

SharedReg849_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg900_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg812_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg812_out;
SharedReg133_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg133_out;
SharedReg739_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg739_out;
SharedReg163_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg163_out;
   MUX_Product37_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg812_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg133_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg739_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg163_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_0_impl_0_out);

   Delay1No376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_0_impl_0_out,
                 Y => Delay1No376_out);

SharedReg943_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg943_out;
SharedReg162_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg162_out;
SharedReg934_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product37_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg943_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg162_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_0_impl_1_out);

   Delay1No377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_0_impl_1_out,
                 Y => Delay1No377_out);

Delay1No378_out_to_Product37_1_impl_parent_implementedSystem_port_0_cast <= Delay1No378_out;
Delay1No379_out_to_Product37_1_impl_parent_implementedSystem_port_1_cast <= Delay1No379_out;
   Product37_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_1_impl_out,
                 X => Delay1No378_out_to_Product37_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No379_out_to_Product37_1_impl_parent_implementedSystem_port_1_cast);

SharedReg166_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg166_out;
SharedReg851_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg851_out;
SharedReg900_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg815_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg815_out;
SharedReg136_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg136_out;
SharedReg722_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg722_out;
   MUX_Product37_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg166_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg851_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg815_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg136_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg722_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_1_impl_0_out);

   Delay1No378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_1_impl_0_out,
                 Y => Delay1No378_out);

SharedReg918_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg943_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg165_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg165_out;
SharedReg934_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product37_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg165_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_1_impl_1_out);

   Delay1No379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_1_impl_1_out,
                 Y => Delay1No379_out);

Delay1No380_out_to_Product37_2_impl_parent_implementedSystem_port_0_cast <= Delay1No380_out;
Delay1No381_out_to_Product37_2_impl_parent_implementedSystem_port_1_cast <= Delay1No381_out;
   Product37_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_2_impl_out,
                 X => Delay1No380_out_to_Product37_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No381_out_to_Product37_2_impl_parent_implementedSystem_port_1_cast);

SharedReg746_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg746_out;
SharedReg169_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg169_out;
SharedReg853_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg853_out;
SharedReg900_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg890_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg890_out;
SharedReg139_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg139_out;
   MUX_Product37_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg746_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg169_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg853_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg890_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg139_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_2_impl_0_out);

   Delay1No380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_2_impl_0_out,
                 Y => Delay1No380_out);

SharedReg913_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg943_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg178_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg934_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product37_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg943_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_2_impl_1_out);

   Delay1No381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_2_impl_1_out,
                 Y => Delay1No381_out);

Delay1No382_out_to_Product37_3_impl_parent_implementedSystem_port_0_cast <= Delay1No382_out;
Delay1No383_out_to_Product37_3_impl_parent_implementedSystem_port_1_cast <= Delay1No383_out;
   Product37_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_3_impl_out,
                 X => Delay1No382_out_to_Product37_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No383_out_to_Product37_3_impl_parent_implementedSystem_port_1_cast);

SharedReg142_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg805_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg805_out;
SharedReg144_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg144_out;
SharedReg840_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg840_out;
SharedReg900_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg882_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg882_out;
   MUX_Product37_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg805_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg144_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg840_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg882_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_3_impl_0_out);

   Delay1No382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_3_impl_0_out,
                 Y => Delay1No382_out);

SharedReg912_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg943_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg180_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg180_out;
SharedReg934_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product37_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg180_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_3_impl_1_out);

   Delay1No383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_3_impl_1_out,
                 Y => Delay1No383_out);

Delay1No384_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast <= Delay1No384_out;
Delay1No385_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast <= Delay1No385_out;
   Product37_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_4_impl_out,
                 X => Delay1No384_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No385_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg825_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg825_out;
SharedReg145_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg145_out;
SharedReg863_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg863_out;
SharedReg132_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg132_out;
SharedReg856_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg856_out;
   MUX_Product37_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg825_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg145_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg863_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg132_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg856_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_4_impl_0_out);

   Delay1No384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_4_impl_0_out,
                 Y => Delay1No384_out);

SharedReg131_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg934_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg913_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg918_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg943_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg943_out;
   MUX_Product37_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg943_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product37_4_impl_1_out);

   Delay1No385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_4_impl_1_out,
                 Y => Delay1No385_out);

Delay1No386_out_to_Subtract8_4_impl_parent_implementedSystem_port_0_cast <= Delay1No386_out;
Delay1No387_out_to_Subtract8_4_impl_parent_implementedSystem_port_1_cast <= Delay1No387_out;
   Subtract8_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_4_impl_out,
                 X => Delay1No386_out_to_Subtract8_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No387_out_to_Subtract8_4_impl_parent_implementedSystem_port_1_cast);

SharedReg315_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg315_out;
SharedReg309_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg309_out;
SharedReg284_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg284_out;
SharedReg653_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg653_out;
SharedReg15_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg309_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg309_out;
   MUX_Subtract8_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg315_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg309_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg284_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg653_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg15_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg309_out_to_MUX_Subtract8_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract8_4_impl_0_out);

   Delay1No386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_4_impl_0_out,
                 Y => Delay1No386_out);

SharedReg349_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg300_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg181_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg181_out;
SharedReg521_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg521_out;
SharedReg31_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg31_out;
Delay3No39_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_6_cast <= Delay3No39_out;
   MUX_Subtract8_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg181_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg521_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg31_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No39_out_to_MUX_Subtract8_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract8_4_impl_1_out);

   Delay1No387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_4_impl_1_out,
                 Y => Delay1No387_out);

Delay1No388_out_to_Add50_4_impl_parent_implementedSystem_port_0_cast <= Delay1No388_out;
Delay1No389_out_to_Add50_4_impl_parent_implementedSystem_port_1_cast <= Delay1No389_out;
   Add50_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add50_4_impl_out,
                 X => Delay1No388_out_to_Add50_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No389_out_to_Add50_4_impl_parent_implementedSystem_port_1_cast);

SharedReg339_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg339_out;
SharedReg705_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg705_out;
SharedReg671_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg671_out;
SharedReg498_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg498_out;
SharedReg518_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg518_out;
SharedReg583_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg583_out;
   MUX_Add50_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg339_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg705_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg671_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg498_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg518_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg583_out_to_MUX_Add50_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add50_4_impl_0_out);

   Delay1No388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add50_4_impl_0_out,
                 Y => Delay1No388_out);

SharedReg344_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg593_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg593_out;
SharedReg715_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg715_out;
SharedReg508_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg508_out;
SharedReg558_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg558_out;
SharedReg714_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg714_out;
   MUX_Add50_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg593_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg715_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg508_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg558_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg714_out_to_MUX_Add50_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add50_4_impl_1_out);

   Delay1No389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add50_4_impl_1_out,
                 Y => Delay1No389_out);

Delay1No390_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No390_out;
Delay1No391_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No391_out;
   Product18_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_0_impl_out,
                 X => Delay1No390_out_to_Product18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No391_out_to_Product18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg947_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg947_out;
SharedReg910_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg920_out;
SharedReg903_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg947_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg920_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_0_impl_0_out);

   Delay1No390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_0_impl_0_out,
                 Y => Delay1No390_out);

SharedReg893_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg893_out;
SharedReg134_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg134_out;
SharedReg120_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg120_out;
SharedReg798_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg798_out;
SharedReg33_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg32_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
   MUX_Product18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg893_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg120_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg798_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg33_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_0_impl_1_out);

   Delay1No391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_0_impl_1_out,
                 Y => Delay1No391_out);

Delay1No392_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No392_out;
Delay1No393_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No393_out;
   Product18_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_1_impl_out,
                 X => Delay1No392_out_to_Product18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No393_out_to_Product18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg947_out;
SharedReg910_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg920_out;
SharedReg903_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg947_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg920_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_1_impl_0_out);

   Delay1No392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_1_impl_0_out,
                 Y => Delay1No392_out);

SharedReg35_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg693_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg693_out;
SharedReg159_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg159_out;
SharedReg137_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg137_out;
SharedReg742_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg742_out;
SharedReg87_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg87_out;
   MUX_Product18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg693_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg159_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg137_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg742_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg87_out_to_MUX_Product18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_1_impl_1_out);

   Delay1No393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_1_impl_1_out,
                 Y => Delay1No393_out);

Delay1No394_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No394_out;
Delay1No395_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No395_out;
   Product18_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_2_impl_out,
                 X => Delay1No394_out_to_Product18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No395_out_to_Product18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg947_out;
SharedReg910_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg920_out;
   MUX_Product18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg947_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg920_out_to_MUX_Product18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_2_impl_0_out);

   Delay1No394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_2_impl_0_out,
                 Y => Delay1No394_out);

SharedReg91_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg38_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg520_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg520_out;
SharedReg168_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
SharedReg126_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg126_out;
SharedReg803_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg803_out;
   MUX_Product18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg520_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg126_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg803_out_to_MUX_Product18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_2_impl_1_out);

   Delay1No395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_2_impl_1_out,
                 Y => Delay1No395_out);

Delay1No396_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast <= Delay1No396_out;
Delay1No397_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast <= Delay1No397_out;
   Product18_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_3_impl_out,
                 X => Delay1No396_out_to_Product18_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No397_out_to_Product18_3_impl_parent_implementedSystem_port_1_cast);

SharedReg920_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg920_out;
SharedReg903_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg947_out;
SharedReg910_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product18_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg920_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg947_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product18_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_3_impl_0_out);

   Delay1No396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_3_impl_0_out,
                 Y => Delay1No396_out);

SharedReg847_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg847_out;
SharedReg42_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg57_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg855_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg143_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg143_out;
SharedReg115_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg115_out;
   MUX_Product18_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg847_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg143_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg115_out_to_MUX_Product18_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_3_impl_1_out);

   Delay1No397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_3_impl_1_out,
                 Y => Delay1No397_out);

Delay1No398_out_to_Product18_4_impl_parent_implementedSystem_port_0_cast <= Delay1No398_out;
Delay1No399_out_to_Product18_4_impl_parent_implementedSystem_port_1_cast <= Delay1No399_out;
   Product18_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product18_4_impl_out,
                 X => Delay1No398_out_to_Product18_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No399_out_to_Product18_4_impl_parent_implementedSystem_port_1_cast);

SharedReg910_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg903_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg908_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg947_out;
   MUX_Product18_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg947_out_to_MUX_Product18_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_4_impl_0_out);

   Delay1No398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_4_impl_0_out,
                 Y => Delay1No398_out);

SharedReg117_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg104_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg104_out;
SharedReg873_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg873_out;
SharedReg73_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg73_out;
SharedReg45_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg45_out;
SharedReg895_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg895_out;
   MUX_Product18_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg873_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg73_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg45_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg895_out_to_MUX_Product18_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product18_4_impl_1_out);

   Delay1No399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product18_4_impl_1_out,
                 Y => Delay1No399_out);

Delay1No400_out_to_Product19_0_impl_parent_implementedSystem_port_0_cast <= Delay1No400_out;
Delay1No401_out_to_Product19_0_impl_parent_implementedSystem_port_1_cast <= Delay1No401_out;
   Product19_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_0_impl_out,
                 X => Delay1No400_out_to_Product19_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No401_out_to_Product19_0_impl_parent_implementedSystem_port_1_cast);

SharedReg947_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg947_out;
SharedReg162_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg162_out;
SharedReg906_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg920_out;
SharedReg913_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg908_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product19_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg947_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg162_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg920_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product19_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_0_impl_0_out);

   Delay1No400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_0_impl_0_out,
                 Y => Delay1No400_out);

SharedReg354_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg354_out;
SharedReg910_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg134_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg134_out;
SharedReg865_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg865_out;
SharedReg33_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg33_out;
SharedReg107_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg107_out;
   MUX_Product19_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg354_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg134_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg865_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg33_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg107_out_to_MUX_Product19_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_0_impl_1_out);

   Delay1No401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_0_impl_1_out,
                 Y => Delay1No401_out);

Delay1No402_out_to_Product19_1_impl_parent_implementedSystem_port_0_cast <= Delay1No402_out;
Delay1No403_out_to_Product19_1_impl_parent_implementedSystem_port_1_cast <= Delay1No403_out;
   Product19_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_1_impl_out,
                 X => Delay1No402_out_to_Product19_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No403_out_to_Product19_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg947_out;
SharedReg165_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg165_out;
SharedReg906_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg920_out;
SharedReg913_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product19_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg947_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg165_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg920_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product19_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_1_impl_0_out);

   Delay1No402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_1_impl_0_out,
                 Y => Delay1No402_out);

SharedReg123_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg357_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg910_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg159_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg159_out;
SharedReg801_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg801_out;
SharedReg87_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg87_out;
   MUX_Product19_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg801_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg87_out_to_MUX_Product19_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_1_impl_1_out);

   Delay1No403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_1_impl_1_out,
                 Y => Delay1No403_out);

Delay1No404_out_to_Product19_2_impl_parent_implementedSystem_port_0_cast <= Delay1No404_out;
Delay1No405_out_to_Product19_2_impl_parent_implementedSystem_port_1_cast <= Delay1No405_out;
   Product19_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_2_impl_out,
                 X => Delay1No404_out_to_Product19_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No405_out_to_Product19_2_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg908_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg947_out;
SharedReg178_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg906_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg920_out;
   MUX_Product19_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg947_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg920_out_to_MUX_Product19_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_2_impl_0_out);

   Delay1No404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_2_impl_0_out,
                 Y => Delay1No404_out);

SharedReg91_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg126_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg126_out;
SharedReg360_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg360_out;
SharedReg910_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg140_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg140_out;
SharedReg858_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg858_out;
   MUX_Product19_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg360_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg858_out_to_MUX_Product19_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_2_impl_1_out);

   Delay1No405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_2_impl_1_out,
                 Y => Delay1No405_out);

Delay1No406_out_to_Product19_3_impl_parent_implementedSystem_port_0_cast <= Delay1No406_out;
Delay1No407_out_to_Product19_3_impl_parent_implementedSystem_port_1_cast <= Delay1No407_out;
   Product19_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_3_impl_out,
                 X => Delay1No406_out_to_Product19_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No407_out_to_Product19_3_impl_parent_implementedSystem_port_1_cast);

SharedReg920_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg920_out;
SharedReg913_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg908_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg947_out;
SharedReg180_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg180_out;
SharedReg906_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product19_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg920_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg947_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg180_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product19_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_3_impl_0_out);

   Delay1No406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_3_impl_0_out,
                 Y => Delay1No406_out);

SharedReg860_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg860_out;
SharedReg42_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg128_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg473_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg473_out;
SharedReg910_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg128_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg128_out;
   MUX_Product19_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg860_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg128_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg473_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg128_out_to_MUX_Product19_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_3_impl_1_out);

   Delay1No407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_3_impl_1_out,
                 Y => Delay1No407_out);

Delay1No408_out_to_Product19_4_impl_parent_implementedSystem_port_0_cast <= Delay1No408_out;
Delay1No409_out_to_Product19_4_impl_parent_implementedSystem_port_1_cast <= Delay1No409_out;
   Product19_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product19_4_impl_out,
                 X => Delay1No408_out_to_Product19_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No409_out_to_Product19_4_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg906_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg920_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg913_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg908_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg947_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg947_out;
   MUX_Product19_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg947_out_to_MUX_Product19_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_4_impl_0_out);

   Delay1No408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_4_impl_0_out,
                 Y => Delay1No408_out);

SharedReg910_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg117_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg883_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg883_out;
SharedReg73_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg73_out;
SharedReg104_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg104_out;
SharedReg897_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg897_out;
   MUX_Product19_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg883_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg73_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg897_out_to_MUX_Product19_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product19_4_impl_1_out);

   Delay1No409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product19_4_impl_1_out,
                 Y => Delay1No409_out);

Delay1No410_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast <= Delay1No410_out;
Delay1No411_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast <= Delay1No411_out;
   Product28_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_0_impl_out,
                 X => Delay1No410_out_to_Product28_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No411_out_to_Product28_0_impl_parent_implementedSystem_port_1_cast);

SharedReg948_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg948_out;
SharedReg900_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg916_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg922_out;
SharedReg903_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg918_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product28_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg948_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg922_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product28_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_0_impl_0_out);

   Delay1No410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_0_impl_0_out,
                 Y => Delay1No410_out);

SharedReg893_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg893_out;
SharedReg172_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg172_out;
SharedReg120_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg120_out;
SharedReg798_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg798_out;
SharedReg812_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg812_out;
SharedReg32_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
   MUX_Product28_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg893_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg172_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg120_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg798_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg812_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product28_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_0_impl_1_out);

   Delay1No411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_0_impl_1_out,
                 Y => Delay1No411_out);

Delay1No412_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast <= Delay1No412_out;
Delay1No413_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast <= Delay1No413_out;
   Product28_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_1_impl_out,
                 X => Delay1No412_out_to_Product28_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No413_out_to_Product28_1_impl_parent_implementedSystem_port_1_cast);

SharedReg918_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg948_out;
SharedReg900_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg916_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg922_out;
SharedReg903_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg903_out;
   MUX_Product28_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg948_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg922_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg903_out_to_MUX_Product28_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_1_impl_0_out);

   Delay1No412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_1_impl_0_out,
                 Y => Delay1No412_out);

SharedReg35_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg693_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg693_out;
SharedReg175_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg175_out;
SharedReg137_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg137_out;
SharedReg742_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg742_out;
SharedReg888_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg888_out;
   MUX_Product28_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg693_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg175_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg137_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg742_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg888_out_to_MUX_Product28_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_1_impl_1_out);

   Delay1No413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_1_impl_1_out,
                 Y => Delay1No413_out);

Delay1No414_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast <= Delay1No414_out;
Delay1No415_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast <= Delay1No415_out;
   Product28_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_2_impl_out,
                 X => Delay1No414_out_to_Product28_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No415_out_to_Product28_2_impl_parent_implementedSystem_port_1_cast);

SharedReg903_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg903_out;
SharedReg918_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg948_out;
SharedReg900_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg916_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg922_out;
   MUX_Product28_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg903_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg948_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg922_out_to_MUX_Product28_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_2_impl_0_out);

   Delay1No414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_2_impl_0_out,
                 Y => Delay1No414_out);

SharedReg890_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg890_out;
SharedReg38_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg520_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg520_out;
SharedReg196_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg196_out;
SharedReg126_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg126_out;
SharedReg803_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg803_out;
   MUX_Product28_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg890_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg520_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg196_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg126_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg803_out_to_MUX_Product28_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_2_impl_1_out);

   Delay1No415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_2_impl_1_out,
                 Y => Delay1No415_out);

Delay1No416_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast <= Delay1No416_out;
Delay1No417_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast <= Delay1No417_out;
   Product28_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_3_impl_out,
                 X => Delay1No416_out_to_Product28_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No417_out_to_Product28_3_impl_parent_implementedSystem_port_1_cast);

SharedReg922_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg922_out;
SharedReg903_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg903_out;
SharedReg918_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg948_out;
SharedReg900_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg916_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product28_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg922_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg903_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg948_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product28_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_3_impl_0_out);

   Delay1No416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_3_impl_0_out,
                 Y => Delay1No416_out);

SharedReg847_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg847_out;
SharedReg892_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg892_out;
SharedReg57_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg855_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg183_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg183_out;
SharedReg115_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg115_out;
   MUX_Product28_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg847_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg892_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg183_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg115_out_to_MUX_Product28_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_3_impl_1_out);

   Delay1No417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_3_impl_1_out,
                 Y => Delay1No417_out);

Delay1No418_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast <= Delay1No418_out;
Delay1No419_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast <= Delay1No419_out;
   Product28_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product28_4_impl_out,
                 X => Delay1No418_out_to_Product28_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No419_out_to_Product28_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg916_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg922_out;
SharedReg903_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg903_out;
SharedReg918_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg948_out;
   MUX_Product28_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg922_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg903_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg948_out_to_MUX_Product28_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_4_impl_0_out);

   Delay1No418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_4_impl_0_out,
                 Y => Delay1No418_out);

SharedReg146_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg146_out;
SharedReg104_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg104_out;
SharedReg873_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg873_out;
SharedReg857_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg857_out;
SharedReg45_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg45_out;
SharedReg895_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg895_out;
   MUX_Product28_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg146_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg873_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg857_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg45_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg895_out_to_MUX_Product28_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product28_4_impl_1_out);

   Delay1No419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product28_4_impl_1_out,
                 Y => Delay1No419_out);

Delay1No420_out_to_Product38_0_impl_parent_implementedSystem_port_0_cast <= Delay1No420_out;
Delay1No421_out_to_Product38_0_impl_parent_implementedSystem_port_1_cast <= Delay1No421_out;
   Product38_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_0_impl_out,
                 X => Delay1No420_out_to_Product38_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No421_out_to_Product38_0_impl_parent_implementedSystem_port_1_cast);

SharedReg354_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg354_out;
SharedReg900_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg134_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg134_out;
SharedReg865_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg865_out;
SharedReg913_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg913_out;
SharedReg107_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg107_out;
   MUX_Product38_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg354_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg134_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg865_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg913_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg107_out_to_MUX_Product38_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_0_impl_0_out);

   Delay1No420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_0_impl_0_out,
                 Y => Delay1No420_out);

SharedReg948_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg948_out;
SharedReg189_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg189_out;
SharedReg916_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg922_out;
SharedReg812_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg812_out;
SharedReg918_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product38_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg948_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg922_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg812_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product38_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_0_impl_1_out);

   Delay1No421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_0_impl_1_out,
                 Y => Delay1No421_out);

Delay1No422_out_to_Product38_1_impl_parent_implementedSystem_port_0_cast <= Delay1No422_out;
Delay1No423_out_to_Product38_1_impl_parent_implementedSystem_port_1_cast <= Delay1No423_out;
   Product38_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_1_impl_out,
                 X => Delay1No422_out_to_Product38_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No423_out_to_Product38_1_impl_parent_implementedSystem_port_1_cast);

SharedReg123_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg123_out;
SharedReg357_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg900_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg159_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg159_out;
SharedReg801_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg801_out;
SharedReg913_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg913_out;
   MUX_Product38_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg123_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg801_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg913_out_to_MUX_Product38_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_1_impl_0_out);

   Delay1No422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_1_impl_0_out,
                 Y => Delay1No422_out);

SharedReg918_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg948_out;
SharedReg200_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg200_out;
SharedReg916_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg922_out;
SharedReg888_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg888_out;
   MUX_Product38_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg948_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg200_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg922_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg888_out_to_MUX_Product38_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_1_impl_1_out);

   Delay1No423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_1_impl_1_out,
                 Y => Delay1No423_out);

Delay1No424_out_to_Product38_2_impl_parent_implementedSystem_port_0_cast <= Delay1No424_out;
Delay1No425_out_to_Product38_2_impl_parent_implementedSystem_port_1_cast <= Delay1No425_out;
   Product38_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_2_impl_out,
                 X => Delay1No424_out_to_Product38_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No425_out_to_Product38_2_impl_parent_implementedSystem_port_1_cast);

SharedReg913_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg913_out;
SharedReg126_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg126_out;
SharedReg360_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg360_out;
SharedReg900_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg140_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg140_out;
SharedReg858_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg858_out;
   MUX_Product38_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg913_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg360_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg140_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg858_out_to_MUX_Product38_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_2_impl_0_out);

   Delay1No424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_2_impl_0_out,
                 Y => Delay1No424_out);

SharedReg890_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg890_out;
SharedReg918_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg948_out;
SharedReg203_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg203_out;
SharedReg916_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg922_out;
   MUX_Product38_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg890_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg948_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg203_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg922_out_to_MUX_Product38_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_2_impl_1_out);

   Delay1No425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_2_impl_1_out,
                 Y => Delay1No425_out);

Delay1No426_out_to_Product38_3_impl_parent_implementedSystem_port_0_cast <= Delay1No426_out;
Delay1No427_out_to_Product38_3_impl_parent_implementedSystem_port_1_cast <= Delay1No427_out;
   Product38_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_3_impl_out,
                 X => Delay1No426_out_to_Product38_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No427_out_to_Product38_3_impl_parent_implementedSystem_port_1_cast);

SharedReg860_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg860_out;
SharedReg913_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg913_out;
SharedReg128_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg473_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg473_out;
SharedReg900_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg128_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg128_out;
   MUX_Product38_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg860_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg913_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg128_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg473_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg128_out_to_MUX_Product38_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_3_impl_0_out);

   Delay1No426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_3_impl_0_out,
                 Y => Delay1No426_out);

SharedReg922_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg922_out;
SharedReg892_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg892_out;
SharedReg918_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg948_out;
SharedReg206_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg916_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product38_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg922_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg892_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg948_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product38_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_3_impl_1_out);

   Delay1No427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_3_impl_1_out,
                 Y => Delay1No427_out);

Delay1No428_out_to_Product38_4_impl_parent_implementedSystem_port_0_cast <= Delay1No428_out;
Delay1No429_out_to_Product38_4_impl_parent_implementedSystem_port_1_cast <= Delay1No429_out;
   Product38_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product38_4_impl_out,
                 X => Delay1No428_out_to_Product38_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No429_out_to_Product38_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg117_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg883_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg883_out;
SharedReg913_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg913_out;
SharedReg104_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg104_out;
SharedReg897_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg897_out;
   MUX_Product38_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg883_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg913_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg897_out_to_MUX_Product38_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_4_impl_0_out);

   Delay1No428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_4_impl_0_out,
                 Y => Delay1No428_out);

SharedReg186_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg916_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg922_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg922_out;
SharedReg857_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg857_out;
SharedReg918_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg948_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg948_out;
   MUX_Product38_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg922_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg857_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg948_out_to_MUX_Product38_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product38_4_impl_1_out);

   Delay1No429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product38_4_impl_1_out,
                 Y => Delay1No429_out);

Delay1No430_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No430_out;
Delay1No431_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No431_out;
   Subtract10_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_3_impl_out,
                 X => Delay1No430_out_to_Subtract10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No431_out_to_Subtract10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg343_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg343_out;
SharedReg265_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg265_out;
SharedReg649_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg649_out;
SharedReg14_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
SharedReg251_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg251_out;
SharedReg307_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg307_out;
   MUX_Subtract10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg343_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg265_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg649_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg14_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg251_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg307_out_to_MUX_Subtract10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract10_3_impl_0_out);

   Delay1No430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_3_impl_0_out,
                 Y => Delay1No430_out);

SharedReg567_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg567_out;
SharedReg170_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg170_out;
SharedReg695_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg695_out;
SharedReg30_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg30_out;
SharedReg154_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg154_out;
SharedReg298_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg298_out;
   MUX_Subtract10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg567_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg695_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg30_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg154_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg298_out_to_MUX_Subtract10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract10_3_impl_1_out);

   Delay1No431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_3_impl_1_out,
                 Y => Delay1No431_out);

Delay1No432_out_to_Add52_0_impl_parent_implementedSystem_port_0_cast <= Delay1No432_out;
Delay1No433_out_to_Add52_0_impl_parent_implementedSystem_port_1_cast <= Delay1No433_out;
   Add52_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add52_0_impl_out,
                 X => Delay1No432_out_to_Add52_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No433_out_to_Add52_0_impl_parent_implementedSystem_port_1_cast);

SharedReg571_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg571_out;
SharedReg335_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg335_out;
SharedReg697_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg697_out;
SharedReg758_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg758_out;
SharedReg688_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg688_out;
SharedReg688_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg688_out;
   MUX_Add52_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg335_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg697_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg758_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg688_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg688_out_to_MUX_Add52_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_0_impl_0_out);

   Delay1No432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_0_impl_0_out,
                 Y => Delay1No432_out);

SharedReg706_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg706_out;
SharedReg340_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg340_out;
SharedReg585_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg585_out;
SharedReg769_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg769_out;
SharedReg696_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg696_out;
SharedReg696_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg696_out;
   MUX_Add52_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg706_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg585_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg769_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg696_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg696_out_to_MUX_Add52_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_0_impl_1_out);

   Delay1No433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_0_impl_1_out,
                 Y => Delay1No433_out);

Delay1No434_out_to_Add52_1_impl_parent_implementedSystem_port_0_cast <= Delay1No434_out;
Delay1No435_out_to_Add52_1_impl_parent_implementedSystem_port_1_cast <= Delay1No435_out;
   Add52_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add52_1_impl_out,
                 X => Delay1No434_out_to_Add52_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No435_out_to_Add52_1_impl_parent_implementedSystem_port_1_cast);

SharedReg689_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg689_out;
SharedReg574_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg574_out;
SharedReg336_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg336_out;
SharedReg699_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg699_out;
SharedReg426_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg426_out;
SharedReg770_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg770_out;
   MUX_Add52_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg689_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg574_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg336_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg699_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg426_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_Add52_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_1_impl_0_out);

   Delay1No434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_1_impl_0_out,
                 Y => Delay1No434_out);

SharedReg698_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg698_out;
SharedReg708_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg708_out;
SharedReg341_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg341_out;
SharedReg587_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg587_out;
SharedReg455_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg455_out;
SharedReg780_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg780_out;
   MUX_Add52_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg698_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg708_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg341_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg587_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg455_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg780_out_to_MUX_Add52_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_1_impl_1_out);

   Delay1No435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_1_impl_1_out,
                 Y => Delay1No435_out);

Delay1No436_out_to_Add52_2_impl_parent_implementedSystem_port_0_cast <= Delay1No436_out;
Delay1No437_out_to_Add52_2_impl_parent_implementedSystem_port_1_cast <= Delay1No437_out;
   Add52_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add52_2_impl_out,
                 X => Delay1No436_out_to_Add52_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No437_out_to_Add52_2_impl_parent_implementedSystem_port_1_cast);

SharedReg772_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg772_out;
SharedReg690_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg690_out;
SharedReg577_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg577_out;
SharedReg337_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg337_out;
SharedReg677_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg677_out;
SharedReg783_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg783_out;
   MUX_Add52_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg772_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg690_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg577_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg337_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg677_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg783_out_to_MUX_Add52_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_2_impl_0_out);

   Delay1No436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_2_impl_0_out,
                 Y => Delay1No436_out);

SharedReg782_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg782_out;
SharedReg700_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg700_out;
SharedReg710_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg710_out;
SharedReg342_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg342_out;
SharedReg685_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg685_out;
SharedReg792_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg792_out;
   MUX_Add52_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg782_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg700_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg710_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg342_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg685_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg792_out_to_MUX_Add52_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_2_impl_1_out);

   Delay1No437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_2_impl_1_out,
                 Y => Delay1No437_out);

Delay1No438_out_to_Add52_3_impl_parent_implementedSystem_port_0_cast <= Delay1No438_out;
Delay1No439_out_to_Add52_3_impl_parent_implementedSystem_port_1_cast <= Delay1No439_out;
   Add52_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add52_3_impl_out,
                 X => Delay1No438_out_to_Add52_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No439_out_to_Add52_3_impl_parent_implementedSystem_port_1_cast);

SharedReg430_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg430_out;
SharedReg691_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg691_out;
SharedReg516_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg516_out;
SharedReg679_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg679_out;
SharedReg338_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg338_out;
SharedReg679_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg679_out;
   MUX_Add52_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg430_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg691_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg516_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg679_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg338_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg679_out_to_MUX_Add52_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_3_impl_0_out);

   Delay1No438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_3_impl_0_out,
                 Y => Delay1No438_out);

SharedReg459_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg459_out;
SharedReg702_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg702_out;
SharedReg556_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg556_out;
SharedReg686_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg686_out;
SharedReg343_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg343_out;
SharedReg686_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg686_out;
   MUX_Add52_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg459_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg702_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg556_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg686_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg343_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg686_out_to_MUX_Add52_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add52_3_impl_1_out);

   Delay1No439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add52_3_impl_1_out,
                 Y => Delay1No439_out);

Delay1No440_out_to_Add54_0_impl_parent_implementedSystem_port_0_cast <= Delay1No440_out;
Delay1No441_out_to_Add54_0_impl_parent_implementedSystem_port_1_cast <= Delay1No441_out;
   Add54_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add54_0_impl_out,
                 X => Delay1No440_out_to_Add54_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No441_out_to_Add54_0_impl_parent_implementedSystem_port_1_cast);

SharedReg664_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg664_out;
SharedReg368_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg368_out;
SharedReg673_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg673_out;
SharedReg424_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg424_out;
SharedReg768_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg768_out;
SharedReg768_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg768_out;
   MUX_Add54_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg664_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg368_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg673_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg424_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg768_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg768_out_to_MUX_Add54_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add54_0_impl_0_out);

   Delay1No440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_0_impl_0_out,
                 Y => Delay1No440_out);

SharedReg768_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg768_out;
SharedReg373_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg373_out;
SharedReg683_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg683_out;
SharedReg453_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg453_out;
SharedReg778_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg778_out;
SharedReg778_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg778_out;
   MUX_Add54_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg768_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg373_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg683_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg453_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg778_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg778_out_to_MUX_Add54_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add54_0_impl_1_out);

   Delay1No441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_0_impl_1_out,
                 Y => Delay1No441_out);

Delay1No442_out_to_Add54_3_impl_parent_implementedSystem_port_0_cast <= Delay1No442_out;
Delay1No443_out_to_Add54_3_impl_parent_implementedSystem_port_1_cast <= Delay1No443_out;
   Add54_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add54_3_impl_out,
                 X => Delay1No442_out_to_Add54_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No443_out_to_Add54_3_impl_parent_implementedSystem_port_1_cast);

SharedReg785_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg785_out;
SharedReg774_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg774_out;
SharedReg691_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg691_out;
SharedReg580_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg580_out;
SharedReg371_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg371_out;
SharedReg775_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg775_out;
   MUX_Add54_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg785_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg774_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg691_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg580_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg371_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg775_out_to_MUX_Add54_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add54_3_impl_0_out);

   Delay1No442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_3_impl_0_out,
                 Y => Delay1No442_out);

SharedReg794_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg794_out;
SharedReg784_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg784_out;
SharedReg702_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg702_out;
SharedReg712_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg712_out;
SharedReg376_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg376_out;
SharedReg785_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg785_out;
   MUX_Add54_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg794_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg784_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg702_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg712_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg376_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg785_out_to_MUX_Add54_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add54_3_impl_1_out);

   Delay1No443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_3_impl_1_out,
                 Y => Delay1No443_out);

Delay1No444_out_to_Add54_4_impl_parent_implementedSystem_port_0_cast <= Delay1No444_out;
Delay1No445_out_to_Add54_4_impl_parent_implementedSystem_port_1_cast <= Delay1No445_out;
   Add54_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add54_4_impl_out,
                 X => Delay1No444_out_to_Add54_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No445_out_to_Add54_4_impl_parent_implementedSystem_port_1_cast);

SharedReg372_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg372_out;
SharedReg681_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg681_out;
SharedReg766_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg766_out;
SharedReg568_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg568_out;
SharedReg692_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg692_out;
SharedReg672_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg672_out;
   MUX_Add54_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg372_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg681_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg766_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg568_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg692_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg672_out_to_MUX_Add54_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add54_4_impl_0_out);

   Delay1No444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_4_impl_0_out,
                 Y => Delay1No444_out);

SharedReg377_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg377_out;
SharedReg687_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg687_out;
SharedReg777_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg777_out;
SharedReg582_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg582_out;
SharedReg704_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg704_out;
SharedReg776_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg776_out;
   MUX_Add54_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg377_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg687_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg777_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg582_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg704_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg776_out_to_MUX_Add54_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add54_4_impl_1_out);

   Delay1No445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_4_impl_1_out,
                 Y => Delay1No445_out);

Delay1No446_out_to_Product42_0_impl_parent_implementedSystem_port_0_cast <= Delay1No446_out;
Delay1No447_out_to_Product42_0_impl_parent_implementedSystem_port_1_cast <= Delay1No447_out;
   Product42_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_0_impl_out,
                 X => Delay1No446_out_to_Product42_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No447_out_to_Product42_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg929_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg926_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product42_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg926_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product42_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_0_impl_0_out);

   Delay1No446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_0_impl_0_out,
                 Y => Delay1No446_out);

SharedReg99_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg172_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg172_out;
SharedReg866_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg866_out;
SharedReg49_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg49_out;
SharedReg875_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg875_out;
SharedReg893_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg893_out;
   MUX_Product42_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg172_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg866_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg49_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg875_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg893_out_to_MUX_Product42_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_0_impl_1_out);

   Delay1No447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_0_impl_1_out,
                 Y => Delay1No447_out);

Delay1No448_out_to_Product42_1_impl_parent_implementedSystem_port_0_cast <= Delay1No448_out;
Delay1No449_out_to_Product42_1_impl_parent_implementedSystem_port_1_cast <= Delay1No449_out;
   Product42_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_1_impl_out,
                 X => Delay1No448_out_to_Product42_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No449_out_to_Product42_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg929_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg926_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg926_out;
   MUX_Product42_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg926_out_to_MUX_Product42_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_1_impl_0_out);

   Delay1No448_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_1_impl_0_out,
                 Y => Delay1No448_out);

SharedReg693_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg693_out;
SharedReg109_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg109_out;
SharedReg175_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg175_out;
SharedReg868_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg868_out;
SharedReg35_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg877_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg877_out;
   MUX_Product42_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg693_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg109_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg175_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg868_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg877_out_to_MUX_Product42_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_1_impl_1_out);

   Delay1No449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_1_impl_1_out,
                 Y => Delay1No449_out);

Delay1No450_out_to_Product42_2_impl_parent_implementedSystem_port_0_cast <= Delay1No450_out;
Delay1No451_out_to_Product42_2_impl_parent_implementedSystem_port_1_cast <= Delay1No451_out;
   Product42_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_2_impl_out,
                 X => Delay1No450_out_to_Product42_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No451_out_to_Product42_2_impl_parent_implementedSystem_port_1_cast);

SharedReg926_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg929_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product42_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg926_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product42_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_2_impl_0_out);

   Delay1No450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_2_impl_0_out,
                 Y => Delay1No450_out);

SharedReg879_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg879_out;
SharedReg520_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg520_out;
SharedReg111_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg111_out;
SharedReg196_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg196_out;
SharedReg859_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg859_out;
SharedReg38_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg38_out;
   MUX_Product42_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg879_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg520_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg111_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg196_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg859_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product42_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_2_impl_1_out);

   Delay1No451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_2_impl_1_out,
                 Y => Delay1No451_out);

Delay1No452_out_to_Product42_3_impl_parent_implementedSystem_port_0_cast <= Delay1No452_out;
Delay1No453_out_to_Product42_3_impl_parent_implementedSystem_port_1_cast <= Delay1No453_out;
   Product42_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_3_impl_out,
                 X => Delay1No452_out_to_Product42_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No453_out_to_Product42_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg926_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg910_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg929_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product42_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg926_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product42_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_3_impl_0_out);

   Delay1No452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_3_impl_0_out,
                 Y => Delay1No452_out);

SharedReg57_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg881_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg881_out;
SharedReg473_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg473_out;
SharedReg101_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg183_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg183_out;
SharedReg848_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg848_out;
   MUX_Product42_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg881_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg473_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg183_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg848_out_to_MUX_Product42_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_3_impl_1_out);

   Delay1No453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_3_impl_1_out,
                 Y => Delay1No453_out);

Delay1No454_out_to_Product42_4_impl_parent_implementedSystem_port_0_cast <= Delay1No454_out;
Delay1No455_out_to_Product42_4_impl_parent_implementedSystem_port_1_cast <= Delay1No455_out;
   Product42_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_4_impl_out,
                 X => Delay1No454_out_to_Product42_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No455_out_to_Product42_4_impl_parent_implementedSystem_port_1_cast);

SharedReg910_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg929_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg902_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg926_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product42_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg926_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product42_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_4_impl_0_out);

   Delay1No454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_4_impl_0_out,
                 Y => Delay1No454_out);

SharedReg146_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg146_out;
SharedReg863_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg863_out;
SharedReg83_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg83_out;
SharedReg883_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg895_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg895_out;
SharedReg94_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg94_out;
   MUX_Product42_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg146_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg863_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg83_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg883_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg895_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Product42_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product42_4_impl_1_out);

   Delay1No455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_4_impl_1_out,
                 Y => Delay1No455_out);

Delay1No456_out_to_Product114_0_impl_parent_implementedSystem_port_0_cast <= Delay1No456_out;
Delay1No457_out_to_Product114_0_impl_parent_implementedSystem_port_1_cast <= Delay1No457_out;
   Product114_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_0_impl_out,
                 X => Delay1No456_out_to_Product114_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No457_out_to_Product114_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg189_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg189_out;
SharedReg929_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg49_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg49_out;
SharedReg875_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg875_out;
SharedReg908_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product114_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg49_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg875_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_0_impl_0_out);

   Delay1No456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_0_impl_0_out,
                 Y => Delay1No456_out);

SharedReg106_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg910_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg876_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg876_out;
SharedReg912_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg931_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg622_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg622_out;
   MUX_Product114_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg876_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg622_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_0_impl_1_out);

   Delay1No457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_0_impl_1_out,
                 Y => Delay1No457_out);

Delay1No458_out_to_Product114_1_impl_parent_implementedSystem_port_0_cast <= Delay1No458_out;
Delay1No459_out_to_Product114_1_impl_parent_implementedSystem_port_1_cast <= Delay1No459_out;
   Product114_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_1_impl_out,
                 X => Delay1No458_out_to_Product114_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No459_out_to_Product114_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg200_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg200_out;
SharedReg929_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg35_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg35_out;
SharedReg877_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg877_out;
   MUX_Product114_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg200_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg35_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg877_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_1_impl_0_out);

   Delay1No458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_1_impl_0_out,
                 Y => Delay1No458_out);

SharedReg612_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg612_out;
SharedReg122_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg122_out;
SharedReg910_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg878_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg878_out;
SharedReg912_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg931_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg931_out;
   MUX_Product114_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg612_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg878_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg931_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_1_impl_1_out);

   Delay1No459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_1_impl_1_out,
                 Y => Delay1No459_out);

Delay1No460_out_to_Product114_2_impl_parent_implementedSystem_port_0_cast <= Delay1No460_out;
Delay1No461_out_to_Product114_2_impl_parent_implementedSystem_port_1_cast <= Delay1No461_out;
   Product114_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_2_impl_out,
                 X => Delay1No460_out_to_Product114_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No461_out_to_Product114_2_impl_parent_implementedSystem_port_1_cast);

SharedReg879_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg879_out;
SharedReg908_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg203_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg203_out;
SharedReg929_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg38_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg38_out;
   MUX_Product114_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg879_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg203_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_2_impl_0_out);

   Delay1No460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_2_impl_0_out,
                 Y => Delay1No460_out);

SharedReg931_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg931_out;
SharedReg616_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg616_out;
SharedReg125_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg910_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg870_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg870_out;
SharedReg912_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product114_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg931_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg616_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg125_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg870_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_2_impl_1_out);

   Delay1No461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_2_impl_1_out,
                 Y => Delay1No461_out);

Delay1No462_out_to_Product114_3_impl_parent_implementedSystem_port_0_cast <= Delay1No462_out;
Delay1No463_out_to_Product114_3_impl_parent_implementedSystem_port_1_cast <= Delay1No463_out;
   Product114_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_3_impl_out,
                 X => Delay1No462_out_to_Product114_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No463_out_to_Product114_3_impl_parent_implementedSystem_port_1_cast);

SharedReg57_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg881_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg881_out;
SharedReg908_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg206_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg929_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product114_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg881_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product114_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_3_impl_0_out);

   Delay1No462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_3_impl_0_out,
                 Y => Delay1No462_out);

SharedReg912_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg931_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg619_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg619_out;
SharedReg114_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg910_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg861_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg861_out;
   MUX_Product114_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg619_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg861_out_to_MUX_Product114_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_3_impl_1_out);

   Delay1No463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_3_impl_1_out,
                 Y => Delay1No463_out);

Delay1No464_out_to_Product114_4_impl_parent_implementedSystem_port_0_cast <= Delay1No464_out;
Delay1No465_out_to_Product114_4_impl_parent_implementedSystem_port_1_cast <= Delay1No465_out;
   Product114_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_4_impl_out,
                 X => Delay1No464_out_to_Product114_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No465_out_to_Product114_4_impl_parent_implementedSystem_port_1_cast);

SharedReg186_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg186_out;
SharedReg929_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg83_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg83_out;
SharedReg883_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg883_out;
SharedReg908_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product114_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg186_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg83_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg883_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product114_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_4_impl_0_out);

   Delay1No464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_4_impl_0_out,
                 Y => Delay1No464_out);

SharedReg910_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg874_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg874_out;
SharedReg912_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg931_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg657_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg657_out;
SharedReg96_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg96_out;
   MUX_Product114_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg874_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg657_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg96_out_to_MUX_Product114_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product114_4_impl_1_out);

   Delay1No465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_4_impl_1_out,
                 Y => Delay1No465_out);

Delay1No466_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast <= Delay1No466_out;
Delay1No467_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast <= Delay1No467_out;
   Product213_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_0_impl_out,
                 X => Delay1No466_out_to_Product213_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No467_out_to_Product213_0_impl_parent_implementedSystem_port_1_cast);

SharedReg909_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg905_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg905_out;
SharedReg934_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg902_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg902_out;
SharedReg942_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg942_out;
SharedReg918_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product213_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg905_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg902_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg942_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product213_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_0_impl_0_out);

   Delay1No466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_0_impl_0_out,
                 Y => Delay1No466_out);

SharedReg99_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg171_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg171_out;
SharedReg866_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg866_out;
SharedReg828_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg828_out;
SharedReg621_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg621_out;
SharedReg893_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg893_out;
   MUX_Product213_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg866_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg828_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg621_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg893_out_to_MUX_Product213_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_0_impl_1_out);

   Delay1No467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_0_impl_1_out,
                 Y => Delay1No467_out);

Delay1No468_out_to_Product213_1_impl_parent_implementedSystem_port_0_cast <= Delay1No468_out;
Delay1No469_out_to_Product213_1_impl_parent_implementedSystem_port_1_cast <= Delay1No469_out;
   Product213_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_1_impl_out,
                 X => Delay1No468_out_to_Product213_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No469_out_to_Product213_1_impl_parent_implementedSystem_port_1_cast);

SharedReg918_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg905_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg905_out;
SharedReg934_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg902_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg902_out;
SharedReg942_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg942_out;
   MUX_Product213_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg905_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg902_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg942_out_to_MUX_Product213_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_1_impl_0_out);

   Delay1No468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_1_impl_0_out,
                 Y => Delay1No468_out);

SharedReg693_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg693_out;
SharedReg109_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg109_out;
SharedReg174_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg174_out;
SharedReg868_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg868_out;
SharedReg814_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg814_out;
SharedReg611_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg611_out;
   MUX_Product213_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg693_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg109_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg868_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg814_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg611_out_to_MUX_Product213_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_1_impl_1_out);

   Delay1No469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_1_impl_1_out,
                 Y => Delay1No469_out);

Delay1No470_out_to_Product213_2_impl_parent_implementedSystem_port_0_cast <= Delay1No470_out;
Delay1No471_out_to_Product213_2_impl_parent_implementedSystem_port_1_cast <= Delay1No471_out;
   Product213_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_2_impl_out,
                 X => Delay1No470_out_to_Product213_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No471_out_to_Product213_2_impl_parent_implementedSystem_port_1_cast);

SharedReg942_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg942_out;
SharedReg918_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg905_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg905_out;
SharedReg934_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg902_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg902_out;
   MUX_Product213_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg942_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg905_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg902_out_to_MUX_Product213_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_2_impl_0_out);

   Delay1No470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_2_impl_0_out,
                 Y => Delay1No470_out);

SharedReg629_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg629_out;
SharedReg520_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg520_out;
SharedReg111_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg111_out;
SharedReg177_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg177_out;
SharedReg859_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg859_out;
SharedReg817_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg817_out;
   MUX_Product213_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg629_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg520_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg111_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg177_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg859_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg817_out_to_MUX_Product213_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_2_impl_1_out);

   Delay1No471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_2_impl_1_out,
                 Y => Delay1No471_out);

Delay1No472_out_to_Product213_3_impl_parent_implementedSystem_port_0_cast <= Delay1No472_out;
Delay1No473_out_to_Product213_3_impl_parent_implementedSystem_port_1_cast <= Delay1No473_out;
   Product213_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_3_impl_out,
                 X => Delay1No472_out_to_Product213_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No473_out_to_Product213_3_impl_parent_implementedSystem_port_1_cast);

SharedReg902_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg902_out;
SharedReg942_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg942_out;
SharedReg918_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg905_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg905_out;
SharedReg934_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product213_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg902_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg942_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg905_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product213_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_3_impl_0_out);

   Delay1No472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_3_impl_0_out,
                 Y => Delay1No472_out);

SharedReg820_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg820_out;
SharedReg651_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg651_out;
SharedReg473_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg473_out;
SharedReg101_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg179_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg179_out;
SharedReg848_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg848_out;
   MUX_Product213_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg820_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg651_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg473_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg179_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg848_out_to_MUX_Product213_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_3_impl_1_out);

   Delay1No473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_3_impl_1_out,
                 Y => Delay1No473_out);

Delay1No474_out_to_Product213_4_impl_parent_implementedSystem_port_0_cast <= Delay1No474_out;
Delay1No475_out_to_Product213_4_impl_parent_implementedSystem_port_1_cast <= Delay1No475_out;
   Product213_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_4_impl_out,
                 X => Delay1No474_out_to_Product213_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No475_out_to_Product213_4_impl_parent_implementedSystem_port_1_cast);

SharedReg905_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg905_out;
SharedReg934_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg902_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg902_out;
SharedReg942_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg942_out;
SharedReg918_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product213_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg905_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg902_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg942_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product213_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_4_impl_0_out);

   Delay1No474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_4_impl_0_out,
                 Y => Delay1No474_out);

SharedReg145_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg863_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg863_out;
SharedReg895_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg895_out;
SharedReg735_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg735_out;
SharedReg895_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg895_out;
SharedReg94_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg94_out;
   MUX_Product213_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg863_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg895_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg735_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg895_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg94_out_to_MUX_Product213_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product213_4_impl_1_out);

   Delay1No475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_4_impl_1_out,
                 Y => Delay1No475_out);

Delay1No476_out_to_Product313_0_impl_parent_implementedSystem_port_0_cast <= Delay1No476_out;
Delay1No477_out_to_Product313_0_impl_parent_implementedSystem_port_1_cast <= Delay1No477_out;
   Product313_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_0_impl_out,
                 X => Delay1No476_out_to_Product313_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No477_out_to_Product313_0_impl_parent_implementedSystem_port_1_cast);

SharedReg106_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg171_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg171_out;
SharedReg876_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg876_out;
SharedReg828_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg828_out;
SharedReg946_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg946_out;
SharedReg622_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg622_out;
   MUX_Product313_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg876_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg828_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg946_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg622_out_to_MUX_Product313_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_0_impl_0_out);

   Delay1No476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_0_impl_0_out,
                 Y => Delay1No476_out);

SharedReg909_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg915_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg915_out;
SharedReg934_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg912_out;
SharedReg621_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg621_out;
SharedReg918_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product313_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg915_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg912_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg621_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product313_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_0_impl_1_out);

   Delay1No477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_0_impl_1_out,
                 Y => Delay1No477_out);

Delay1No478_out_to_Product313_1_impl_parent_implementedSystem_port_0_cast <= Delay1No478_out;
Delay1No479_out_to_Product313_1_impl_parent_implementedSystem_port_1_cast <= Delay1No479_out;
   Product313_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_1_impl_out,
                 X => Delay1No478_out_to_Product313_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No479_out_to_Product313_1_impl_parent_implementedSystem_port_1_cast);

SharedReg612_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg612_out;
SharedReg122_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg122_out;
SharedReg174_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
SharedReg878_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg878_out;
SharedReg814_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg814_out;
SharedReg946_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg946_out;
   MUX_Product313_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg612_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg122_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg878_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg814_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg946_out_to_MUX_Product313_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_1_impl_0_out);

   Delay1No478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_1_impl_0_out,
                 Y => Delay1No478_out);

SharedReg918_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg915_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg915_out;
SharedReg934_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg912_out;
SharedReg611_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg611_out;
   MUX_Product313_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg915_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg912_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg611_out_to_MUX_Product313_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_1_impl_1_out);

   Delay1No479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_1_impl_1_out,
                 Y => Delay1No479_out);

Delay1No480_out_to_Product313_2_impl_parent_implementedSystem_port_0_cast <= Delay1No480_out;
Delay1No481_out_to_Product313_2_impl_parent_implementedSystem_port_1_cast <= Delay1No481_out;
   Product313_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_2_impl_out,
                 X => Delay1No480_out_to_Product313_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No481_out_to_Product313_2_impl_parent_implementedSystem_port_1_cast);

SharedReg946_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg946_out;
SharedReg616_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg616_out;
SharedReg125_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg177_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg177_out;
SharedReg870_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg870_out;
SharedReg817_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg817_out;
   MUX_Product313_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg946_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg616_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg125_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg177_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg870_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg817_out_to_MUX_Product313_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_2_impl_0_out);

   Delay1No480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_2_impl_0_out,
                 Y => Delay1No480_out);

SharedReg629_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg629_out;
SharedReg918_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg915_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg915_out;
SharedReg934_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg912_out;
   MUX_Product313_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg629_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg915_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg912_out_to_MUX_Product313_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_2_impl_1_out);

   Delay1No481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_2_impl_1_out,
                 Y => Delay1No481_out);

Delay1No482_out_to_Product313_3_impl_parent_implementedSystem_port_0_cast <= Delay1No482_out;
Delay1No483_out_to_Product313_3_impl_parent_implementedSystem_port_1_cast <= Delay1No483_out;
   Product313_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_3_impl_out,
                 X => Delay1No482_out_to_Product313_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No483_out_to_Product313_3_impl_parent_implementedSystem_port_1_cast);

SharedReg820_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg820_out;
SharedReg946_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg946_out;
SharedReg619_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg619_out;
SharedReg114_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
SharedReg179_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg179_out;
SharedReg861_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg861_out;
   MUX_Product313_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg820_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg946_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg619_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg179_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg861_out_to_MUX_Product313_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_3_impl_0_out);

   Delay1No482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_3_impl_0_out,
                 Y => Delay1No482_out);

SharedReg912_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg912_out;
SharedReg651_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg651_out;
SharedReg918_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg915_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg915_out;
SharedReg934_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product313_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg912_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg651_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg915_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product313_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_3_impl_1_out);

   Delay1No483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_3_impl_1_out,
                 Y => Delay1No483_out);

Delay1No484_out_to_Product313_4_impl_parent_implementedSystem_port_0_cast <= Delay1No484_out;
Delay1No485_out_to_Product313_4_impl_parent_implementedSystem_port_1_cast <= Delay1No485_out;
   Product313_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_4_impl_out,
                 X => Delay1No484_out_to_Product313_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No485_out_to_Product313_4_impl_parent_implementedSystem_port_1_cast);

SharedReg145_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg874_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg874_out;
SharedReg895_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg895_out;
SharedReg946_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg946_out;
SharedReg657_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg657_out;
SharedReg96_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg96_out;
   MUX_Product313_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg874_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg895_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg946_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg657_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg96_out_to_MUX_Product313_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_4_impl_0_out);

   Delay1No484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_4_impl_0_out,
                 Y => Delay1No484_out);

SharedReg915_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg915_out;
SharedReg934_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg912_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg912_out;
SharedReg735_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg735_out;
SharedReg918_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product313_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg915_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg912_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg735_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product313_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product313_4_impl_1_out);

   Delay1No485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_4_impl_1_out,
                 Y => Delay1No485_out);

Delay1No486_out_to_Subtract14_4_impl_parent_implementedSystem_port_0_cast <= Delay1No486_out;
Delay1No487_out_to_Subtract14_4_impl_parent_implementedSystem_port_1_cast <= Delay1No487_out;
   Subtract14_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract14_4_impl_out,
                 X => Delay1No486_out_to_Subtract14_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No487_out_to_Subtract14_4_impl_parent_implementedSystem_port_1_cast);

SharedReg2_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg2_out;
SharedReg489_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg489_out;
SharedReg786_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg786_out;
SharedReg558_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg558_out;
Delay3No149_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_5_cast <= Delay3No149_out;
SharedReg422_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg422_out;
   MUX_Subtract14_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg489_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg786_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg558_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No149_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg422_out_to_MUX_Subtract14_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract14_4_impl_0_out);

   Delay1No486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract14_4_impl_0_out,
                 Y => Delay1No486_out);

SharedReg18_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg519_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg519_out;
SharedReg797_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg797_out;
SharedReg593_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg593_out;
Delay3No154_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_5_cast <= Delay3No154_out;
SharedReg471_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg471_out;
   MUX_Subtract14_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg519_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg797_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg593_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No154_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg471_out_to_MUX_Subtract14_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract14_4_impl_1_out);

   Delay1No487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract14_4_impl_1_out,
                 Y => Delay1No487_out);

Delay1No488_out_to_Subtract17_0_impl_parent_implementedSystem_port_0_cast <= Delay1No488_out;
Delay1No489_out_to_Subtract17_0_impl_parent_implementedSystem_port_1_cast <= Delay1No489_out;
   Subtract17_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract17_0_impl_out,
                 X => Delay1No488_out_to_Subtract17_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No489_out_to_Subtract17_0_impl_parent_implementedSystem_port_1_cast);

Delay4No70_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_1_cast <= Delay4No70_out;
SharedReg1_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg414_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg414_out;
SharedReg778_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg778_out;
SharedReg683_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg683_out;
Delay3No145_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_6_cast <= Delay3No145_out;
   MUX_Subtract17_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No70_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg414_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg778_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg683_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No145_out_to_MUX_Subtract17_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract17_0_impl_0_out);

   Delay1No488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_0_impl_0_out,
                 Y => Delay1No488_out);

Delay4No85_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_1_cast <= Delay4No85_out;
SharedReg17_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg463_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg463_out;
SharedReg789_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg789_out;
SharedReg706_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg706_out;
Delay3No150_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_6_cast <= Delay3No150_out;
   MUX_Subtract17_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No85_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg463_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg789_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg706_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No150_out_to_MUX_Subtract17_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract17_0_impl_1_out);

   Delay1No489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_0_impl_1_out,
                 Y => Delay1No489_out);

Delay1No490_out_to_Subtract17_1_impl_parent_implementedSystem_port_0_cast <= Delay1No490_out;
Delay1No491_out_to_Subtract17_1_impl_parent_implementedSystem_port_1_cast <= Delay1No491_out;
   Subtract17_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract17_1_impl_out,
                 X => Delay1No490_out_to_Subtract17_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No491_out_to_Subtract17_1_impl_parent_implementedSystem_port_1_cast);

Delay3No146_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No146_out;
Delay4No71_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No71_out;
SharedReg1_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg416_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg416_out;
SharedReg201_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg201_out;
SharedReg760_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg760_out;
   MUX_Subtract17_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No146_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No71_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg416_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg201_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg760_out_to_MUX_Subtract17_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract17_1_impl_0_out);

   Delay1No490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_1_impl_0_out,
                 Y => Delay1No490_out);

Delay3No151_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_1_cast <= Delay3No151_out;
Delay4No86_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_2_cast <= Delay4No86_out;
SharedReg17_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
SharedReg465_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg465_out;
SharedReg214_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg214_out;
SharedReg790_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg790_out;
   MUX_Subtract17_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No151_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No86_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg17_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg465_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg214_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg790_out_to_MUX_Subtract17_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract17_1_impl_1_out);

   Delay1No491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract17_1_impl_1_out,
                 Y => Delay1No491_out);

Delay1No492_out_to_Subtract18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No492_out;
Delay1No493_out_to_Subtract18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No493_out;
   Subtract18_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_0_impl_out,
                 X => Delay1No492_out_to_Subtract18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No493_out_to_Subtract18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg414_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg2_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg481_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg481_out;
SharedReg190_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg190_out;
SharedReg758_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg758_out;
SharedReg453_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg453_out;
   MUX_Subtract18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg481_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg190_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg758_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg453_out_to_MUX_Subtract18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract18_0_impl_0_out);

   Delay1No492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_0_impl_0_out,
                 Y => Delay1No492_out);

SharedReg463_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg463_out;
SharedReg18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg511_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg511_out;
SharedReg224_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg224_out;
SharedReg788_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg788_out;
SharedReg490_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg490_out;
   MUX_Subtract18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg463_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg511_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg224_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg788_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg490_out_to_MUX_Subtract18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract18_0_impl_1_out);

   Delay1No493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_0_impl_1_out,
                 Y => Delay1No493_out);

Delay1No494_out_to_Subtract18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No494_out;
Delay1No495_out_to_Subtract18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No495_out;
   Subtract18_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_1_impl_out,
                 X => Delay1No494_out_to_Subtract18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No495_out_to_Subtract18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg455_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg455_out;
SharedReg416_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg416_out;
SharedReg2_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg483_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg483_out;
SharedReg227_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg227_out;
SharedReg610_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg610_out;
   MUX_Subtract18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg455_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg416_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg483_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg227_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg610_out_to_MUX_Subtract18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract18_1_impl_0_out);

   Delay1No494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_1_impl_0_out,
                 Y => Delay1No494_out);

SharedReg492_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg492_out;
SharedReg465_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg465_out;
SharedReg18_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg18_out;
SharedReg513_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg513_out;
SharedReg248_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg248_out;
SharedReg801_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg801_out;
   MUX_Subtract18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg492_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg465_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg18_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg513_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg248_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg801_out_to_MUX_Subtract18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract18_1_impl_1_out);

   Delay1No495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_1_impl_1_out,
                 Y => Delay1No495_out);

Delay1No496_out_to_Subtract18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No496_out;
Delay1No497_out_to_Subtract18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No497_out;
   Subtract18_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract18_2_impl_out,
                 X => Delay1No496_out_to_Subtract18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No497_out_to_Subtract18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg762_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg762_out;
Delay3No147_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_2_cast <= Delay3No147_out;
Delay4No72_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_3_cast <= Delay4No72_out;
SharedReg1_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1_out;
SharedReg485_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg485_out;
SharedReg218_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg218_out;
   MUX_Subtract18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg762_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No147_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No72_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg485_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg218_out_to_MUX_Subtract18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract18_2_impl_0_out);

   Delay1No496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_2_impl_0_out,
                 Y => Delay1No496_out);

SharedReg792_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg792_out;
Delay3No152_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_2_cast <= Delay3No152_out;
Delay4No87_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No87_out;
SharedReg17_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
SharedReg515_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg515_out;
SharedReg232_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg232_out;
   MUX_Subtract18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg792_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No152_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No87_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg515_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg232_out_to_MUX_Subtract18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract18_2_impl_1_out);

   Delay1No497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract18_2_impl_1_out,
                 Y => Delay1No497_out);

Delay1No498_out_to_Subtract19_3_impl_parent_implementedSystem_port_0_cast <= Delay1No498_out;
Delay1No499_out_to_Subtract19_3_impl_parent_implementedSystem_port_1_cast <= Delay1No499_out;
   Subtract19_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract19_3_impl_out,
                 X => Delay1No498_out_to_Subtract19_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No499_out_to_Subtract19_3_impl_parent_implementedSystem_port_1_cast);

SharedReg237_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg237_out;
SharedReg764_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg764_out;
Delay3No148_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_3_cast <= Delay3No148_out;
Delay4No73_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_4_cast <= Delay4No73_out;
SharedReg2_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg486_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg486_out;
   MUX_Subtract19_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg237_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg764_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No148_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No73_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg486_out_to_MUX_Subtract19_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract19_3_impl_0_out);

   Delay1No498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract19_3_impl_0_out,
                 Y => Delay1No498_out);

SharedReg253_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg253_out;
SharedReg794_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg794_out;
Delay3No153_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_3_cast <= Delay3No153_out;
Delay4No88_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_4_cast <= Delay4No88_out;
SharedReg18_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg567_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg567_out;
   MUX_Subtract19_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg253_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg794_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No153_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay4No88_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg567_out_to_MUX_Subtract19_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract19_3_impl_1_out);

   Delay1No499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract19_3_impl_1_out,
                 Y => Delay1No499_out);

Delay1No500_out_to_Subtract20_0_impl_parent_implementedSystem_port_0_cast <= Delay1No500_out;
Delay1No501_out_to_Subtract20_0_impl_parent_implementedSystem_port_1_cast <= Delay1No501_out;
   Subtract20_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_0_impl_out,
                 X => Delay1No500_out_to_Subtract20_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No501_out_to_Subtract20_0_impl_parent_implementedSystem_port_1_cast);

SharedReg480_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg480_out;
SharedReg3_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg480_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg480_out;
SharedReg245_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg245_out;
SharedReg606_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg606_out;
Delay3No195_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_6_cast <= Delay3No195_out;
   MUX_Subtract20_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg480_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg480_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg245_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg606_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No195_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_0_impl_0_out);

   Delay1No500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_0_impl_0_out,
                 Y => Delay1No500_out);

SharedReg510_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg510_out;
SharedReg19_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg561_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg561_out;
SharedReg259_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg259_out;
SharedReg798_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg798_out;
Delay3No210_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_6_cast <= Delay3No210_out;
   MUX_Subtract20_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg510_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg561_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg259_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg798_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No210_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_0_impl_1_out);

   Delay1No501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_0_impl_1_out,
                 Y => Delay1No501_out);

Delay1No502_out_to_Subtract20_1_impl_parent_implementedSystem_port_0_cast <= Delay1No502_out;
Delay1No503_out_to_Subtract20_1_impl_parent_implementedSystem_port_1_cast <= Delay1No503_out;
   Subtract20_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_1_impl_out,
                 X => Delay1No502_out_to_Subtract20_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No503_out_to_Subtract20_1_impl_parent_implementedSystem_port_1_cast);

Delay3No196_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No196_out;
SharedReg482_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg482_out;
SharedReg3_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg482_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg482_out;
SharedReg322_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg322_out;
SharedReg247_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg247_out;
   MUX_Subtract20_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No196_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg482_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg3_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg482_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg322_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg247_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_1_impl_0_out);

   Delay1No502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_1_impl_0_out,
                 Y => Delay1No502_out);

Delay3No211_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_1_cast <= Delay3No211_out;
SharedReg512_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg512_out;
SharedReg19_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg563_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg563_out;
SharedReg407_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg407_out;
SharedReg148_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg148_out;
   MUX_Subtract20_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No211_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg512_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg19_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg563_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg407_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg148_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_1_impl_1_out);

   Delay1No503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_1_impl_1_out,
                 Y => Delay1No503_out);

Delay1No504_out_to_Subtract20_2_impl_parent_implementedSystem_port_0_cast <= Delay1No504_out;
Delay1No505_out_to_Subtract20_2_impl_parent_implementedSystem_port_1_cast <= Delay1No505_out;
   Subtract20_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_2_impl_out,
                 X => Delay1No504_out_to_Subtract20_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No505_out_to_Subtract20_2_impl_parent_implementedSystem_port_1_cast);

SharedReg628_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg628_out;
SharedReg457_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg457_out;
SharedReg418_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg418_out;
SharedReg2_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg2_out;
SharedReg484_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg484_out;
SharedReg389_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg389_out;
   MUX_Subtract20_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg628_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg457_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg418_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg484_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg389_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_2_impl_0_out);

   Delay1No504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_2_impl_0_out,
                 Y => Delay1No504_out);

SharedReg858_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg858_out;
SharedReg494_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg494_out;
SharedReg467_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg467_out;
SharedReg18_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg18_out;
SharedReg565_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg565_out;
SharedReg326_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg326_out;
   MUX_Subtract20_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg858_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg494_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg467_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg18_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg565_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg326_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_2_impl_1_out);

   Delay1No505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_2_impl_1_out,
                 Y => Delay1No505_out);

Delay1No506_out_to_Subtract20_4_impl_parent_implementedSystem_port_0_cast <= Delay1No506_out;
Delay1No507_out_to_Subtract20_4_impl_parent_implementedSystem_port_1_cast <= Delay1No507_out;
   Subtract20_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_4_impl_out,
                 X => Delay1No506_out_to_Subtract20_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No507_out_to_Subtract20_4_impl_parent_implementedSystem_port_1_cast);

SharedReg3_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg488_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg488_out;
SharedReg187_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg187_out;
SharedReg687_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg687_out;
SharedReg461_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg461_out;
SharedReg488_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg488_out;
   MUX_Subtract20_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg488_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg187_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg687_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg461_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg488_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_4_impl_0_out);

   Delay1No506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_4_impl_0_out,
                 Y => Delay1No506_out);

SharedReg19_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg569_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg569_out;
SharedReg258_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg258_out;
SharedReg714_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg714_out;
SharedReg498_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg498_out;
SharedReg518_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg518_out;
   MUX_Subtract20_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg569_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg258_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg714_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg498_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg518_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract20_4_impl_1_out);

   Delay1No507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_4_impl_1_out,
                 Y => Delay1No507_out);

Delay1No508_out_to_Subtract21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No508_out;
Delay1No509_out_to_Subtract21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No509_out;
   Subtract21_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract21_0_impl_out,
                 X => Delay1No508_out_to_Subtract21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No509_out_to_Subtract21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg550_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg550_out;
SharedReg4_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg500_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg500_out;
SharedReg318_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg318_out;
SharedReg244_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg244_out;
SharedReg500_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg500_out;
   MUX_Subtract21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg550_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg500_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg318_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg244_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg500_out_to_MUX_Subtract21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_0_impl_0_out);

   Delay1No508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_0_impl_0_out,
                 Y => Delay1No508_out);

SharedReg585_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg585_out;
SharedReg20_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg586_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg586_out;
SharedReg404_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg404_out;
SharedReg538_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg538_out;
SharedReg560_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg560_out;
   MUX_Subtract21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg585_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg586_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg404_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg538_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg560_out_to_MUX_Subtract21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_0_impl_1_out);

   Delay1No509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_0_impl_1_out,
                 Y => Delay1No509_out);

Delay1No510_out_to_Subtract21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No510_out;
Delay1No511_out_to_Subtract21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No511_out;
   Subtract21_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract21_1_impl_out,
                 X => Delay1No510_out_to_Subtract21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No511_out_to_Subtract21_1_impl_parent_implementedSystem_port_1_cast);

SharedReg502_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg502_out;
SharedReg552_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg552_out;
SharedReg4_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg4_out;
SharedReg502_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg502_out;
SharedReg200_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg200_out;
SharedReg439_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg439_out;
   MUX_Subtract21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg502_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg552_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg4_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg502_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg200_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg439_out_to_MUX_Subtract21_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_1_impl_0_out);

   Delay1No510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_1_impl_0_out,
                 Y => Delay1No510_out);

SharedReg562_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg562_out;
SharedReg587_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg587_out;
SharedReg20_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg588_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg588_out;
SharedReg215_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg215_out;
SharedReg405_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg405_out;
   MUX_Subtract21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg562_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg587_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg588_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg215_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg405_out_to_MUX_Subtract21_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_1_impl_1_out);

   Delay1No511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_1_impl_1_out,
                 Y => Delay1No511_out);

Delay1No512_out_to_Subtract21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No512_out;
Delay1No513_out_to_Subtract21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No513_out;
   Subtract21_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract21_2_impl_out,
                 X => Delay1No512_out_to_Subtract21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No513_out_to_Subtract21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg250_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg250_out;
Delay3No197_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_2_cast <= Delay3No197_out;
SharedReg484_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg484_out;
SharedReg3_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
SharedReg504_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg504_out;
SharedReg196_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg196_out;
   MUX_Subtract21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg250_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No197_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg484_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg3_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg504_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg196_out_to_MUX_Subtract21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_2_impl_0_out);

   Delay1No512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_2_impl_0_out,
                 Y => Delay1No512_out);

SharedReg153_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
Delay3No212_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_2_cast <= Delay3No212_out;
SharedReg514_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg514_out;
SharedReg19_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg19_out;
SharedReg590_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg590_out;
SharedReg204_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg204_out;
   MUX_Subtract21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No212_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg514_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg19_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg590_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg204_out_to_MUX_Subtract21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_2_impl_1_out);

   Delay1No513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_2_impl_1_out,
                 Y => Delay1No513_out);

Delay1No514_out_to_Subtract21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No514_out;
Delay1No515_out_to_Subtract21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No515_out;
   Subtract21_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract21_3_impl_out,
                 X => Delay1No514_out_to_Subtract21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No515_out_to_Subtract21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg362_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg362_out;
SharedReg650_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg650_out;
SharedReg459_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg459_out;
SharedReg420_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg420_out;
SharedReg3_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg506_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg506_out;
   MUX_Subtract21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg362_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg650_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg459_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg420_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg506_out_to_MUX_Subtract21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_3_impl_0_out);

   Delay1No514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_3_impl_0_out,
                 Y => Delay1No514_out);

SharedReg392_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg860_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg860_out;
SharedReg496_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg496_out;
SharedReg469_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg469_out;
SharedReg19_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg19_out;
SharedReg592_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg592_out;
   MUX_Subtract21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg860_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg496_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg469_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg19_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg592_out_to_MUX_Subtract21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_3_impl_1_out);

   Delay1No515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_3_impl_1_out,
                 Y => Delay1No515_out);

Delay1No516_out_to_Subtract21_4_impl_parent_implementedSystem_port_0_cast <= Delay1No516_out;
Delay1No517_out_to_Subtract21_4_impl_parent_implementedSystem_port_1_cast <= Delay1No517_out;
   Subtract21_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract21_4_impl_out,
                 X => Delay1No516_out_to_Subtract21_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No517_out_to_Subtract21_4_impl_parent_implementedSystem_port_1_cast);

SharedReg4_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg508_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg508_out;
SharedReg271_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg271_out;
SharedReg766_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg766_out;
Delay3No199_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_5_cast <= Delay3No199_out;
SharedReg558_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg558_out;
   MUX_Subtract21_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg508_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg271_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg766_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No199_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg558_out_to_MUX_Subtract21_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_4_impl_0_out);

   Delay1No516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_4_impl_0_out,
                 Y => Delay1No516_out);

SharedReg20_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg594_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg594_out;
SharedReg287_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg287_out;
SharedReg796_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg796_out;
Delay3No214_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_5_cast <= Delay3No214_out;
SharedReg593_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg593_out;
   MUX_Subtract21_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg594_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg287_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg796_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No214_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg593_out_to_MUX_Subtract21_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract21_4_impl_1_out);

   Delay1No517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_4_impl_1_out,
                 Y => Delay1No517_out);

Delay1No518_out_to_Add63_4_impl_parent_implementedSystem_port_0_cast <= Delay1No518_out;
Delay1No519_out_to_Add63_4_impl_parent_implementedSystem_port_1_cast <= Delay1No519_out;
   Add63_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add63_4_impl_out,
                 X => Delay1No518_out_to_Add63_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No519_out_to_Add63_4_impl_parent_implementedSystem_port_1_cast);

SharedReg681_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg681_out;
SharedReg777_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg777_out;
SharedReg432_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg432_out;
SharedReg692_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg692_out;
SharedReg776_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg776_out;
Delay3No234_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_6_cast <= Delay3No234_out;
   MUX_Add63_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg681_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg777_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg432_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg692_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg776_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No234_out_to_MUX_Add63_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add63_4_impl_0_out);

   Delay1No518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add63_4_impl_0_out,
                 Y => Delay1No518_out);

SharedReg687_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg687_out;
SharedReg787_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg787_out;
SharedReg461_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg461_out;
SharedReg704_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg704_out;
SharedReg786_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg786_out;
SharedReg796_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg796_out;
   MUX_Add63_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg687_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg787_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg461_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg704_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg786_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg796_out_to_MUX_Add63_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Add63_4_impl_1_out);

   Delay1No519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add63_4_impl_1_out,
                 Y => Delay1No519_out);

Delay1No520_out_to_Product50_0_impl_parent_implementedSystem_port_0_cast <= Delay1No520_out;
Delay1No521_out_to_Product50_0_impl_parent_implementedSystem_port_1_cast <= Delay1No521_out;
   Product50_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_0_impl_out,
                 X => Delay1No520_out_to_Product50_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No521_out_to_Product50_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg928_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg928_out;
SharedReg929_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product50_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg928_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg920_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg926_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product50_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_0_impl_0_out);

   Delay1No520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_0_impl_0_out,
                 Y => Delay1No520_out);

SharedReg244_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg354_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg354_out;
SharedReg829_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg829_out;
SharedReg849_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg849_out;
SharedReg885_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg885_out;
SharedReg51_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg51_out;
   MUX_Product50_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg354_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg829_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg885_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg51_out_to_MUX_Product50_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_0_impl_1_out);

   Delay1No521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_0_impl_1_out,
                 Y => Delay1No521_out);

Delay1No522_out_to_Product50_1_impl_parent_implementedSystem_port_0_cast <= Delay1No522_out;
Delay1No523_out_to_Product50_1_impl_parent_implementedSystem_port_1_cast <= Delay1No523_out;
   Product50_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_1_impl_out,
                 X => Delay1No522_out_to_Product50_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No523_out_to_Product50_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg928_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg928_out;
SharedReg929_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg926_out;
   MUX_Product50_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg928_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg920_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg926_out_to_MUX_Product50_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_1_impl_0_out);

   Delay1No522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_1_impl_0_out,
                 Y => Delay1No522_out);

SharedReg37_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg247_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg247_out;
SharedReg357_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg357_out;
SharedReg833_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg833_out;
SharedReg832_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg832_out;
SharedReg887_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg887_out;
   MUX_Product50_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg247_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg357_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg833_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg832_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg887_out_to_MUX_Product50_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_1_impl_1_out);

   Delay1No523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_1_impl_1_out,
                 Y => Delay1No523_out);

Delay1No524_out_to_Product50_2_impl_parent_implementedSystem_port_0_cast <= Delay1No524_out;
Delay1No525_out_to_Product50_2_impl_parent_implementedSystem_port_1_cast <= Delay1No525_out;
   Product50_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_2_impl_out,
                 X => Delay1No524_out_to_Product50_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No525_out_to_Product50_2_impl_parent_implementedSystem_port_1_cast);

SharedReg926_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg928_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg928_out;
SharedReg929_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg920_out;
   MUX_Product50_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg926_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg928_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg920_out_to_MUX_Product50_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_2_impl_0_out);

   Delay1No524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_2_impl_0_out,
                 Y => Delay1No524_out);

SharedReg889_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg889_out;
SharedReg93_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg93_out;
SharedReg250_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg250_out;
SharedReg520_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg520_out;
SharedReg818_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg818_out;
SharedReg836_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg836_out;
   MUX_Product50_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg889_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg250_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg520_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg818_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg836_out_to_MUX_Product50_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_2_impl_1_out);

   Delay1No525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_2_impl_1_out,
                 Y => Delay1No525_out);

Delay1No526_out_to_Product50_3_impl_parent_implementedSystem_port_0_cast <= Delay1No526_out;
Delay1No527_out_to_Product50_3_impl_parent_implementedSystem_port_1_cast <= Delay1No527_out;
   Product50_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_3_impl_out,
                 X => Delay1No526_out_to_Product50_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No527_out_to_Product50_3_impl_parent_implementedSystem_port_1_cast);

SharedReg920_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg928_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg928_out;
SharedReg929_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product50_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg920_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg926_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg928_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product50_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_3_impl_0_out);

   Delay1No526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_3_impl_0_out,
                 Y => Delay1No526_out);

SharedReg840_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg840_out;
SharedReg891_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg891_out;
SharedReg44_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg44_out;
SharedReg252_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg252_out;
SharedReg855_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg892_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg892_out;
   MUX_Product50_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg840_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg891_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg44_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg892_out_to_MUX_Product50_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_3_impl_1_out);

   Delay1No527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_3_impl_1_out,
                 Y => Delay1No527_out);

Delay1No528_out_to_Product50_4_impl_parent_implementedSystem_port_0_cast <= Delay1No528_out;
Delay1No529_out_to_Product50_4_impl_parent_implementedSystem_port_1_cast <= Delay1No529_out;
   Product50_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product50_4_impl_out,
                 X => Delay1No528_out_to_Product50_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No529_out_to_Product50_4_impl_parent_implementedSystem_port_1_cast);

SharedReg928_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg928_out;
SharedReg929_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg926_out;
SharedReg908_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product50_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg928_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg926_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product50_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_4_impl_0_out);

   Delay1No528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_4_impl_0_out,
                 Y => Delay1No528_out);

SharedReg897_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg897_out;
SharedReg844_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg844_out;
SharedReg897_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg897_out;
SharedReg824_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg824_out;
SharedReg74_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg74_out;
SharedReg257_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg257_out;
   MUX_Product50_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg897_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg844_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg897_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg824_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg74_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg257_out_to_MUX_Product50_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product50_4_impl_1_out);

   Delay1No529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product50_4_impl_1_out,
                 Y => Delay1No529_out);

Delay1No530_out_to_Product122_0_impl_parent_implementedSystem_port_0_cast <= Delay1No530_out;
Delay1No531_out_to_Product122_0_impl_parent_implementedSystem_port_1_cast <= Delay1No531_out;
   Product122_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_0_impl_out,
                 X => Delay1No530_out_to_Product122_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No531_out_to_Product122_0_impl_parent_implementedSystem_port_1_cast);

SharedReg244_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg244_out;
SharedReg354_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg354_out;
SharedReg929_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg926_out;
SharedReg51_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg51_out;
   MUX_Product122_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg244_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg354_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg920_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg926_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg51_out_to_MUX_Product122_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_0_impl_0_out);

   Delay1No530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_0_impl_0_out,
                 Y => Delay1No530_out);

SharedReg909_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg933_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg933_out;
SharedReg850_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg850_out;
SharedReg893_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg893_out;
SharedReg811_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg811_out;
SharedReg918_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product122_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg933_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg850_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg893_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg811_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product122_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_0_impl_1_out);

   Delay1No531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_0_impl_1_out,
                 Y => Delay1No531_out);

Delay1No532_out_to_Product122_1_impl_parent_implementedSystem_port_0_cast <= Delay1No532_out;
Delay1No533_out_to_Product122_1_impl_parent_implementedSystem_port_1_cast <= Delay1No533_out;
   Product122_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_1_impl_out,
                 X => Delay1No532_out_to_Product122_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No533_out_to_Product122_1_impl_parent_implementedSystem_port_1_cast);

SharedReg37_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg247_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg247_out;
SharedReg357_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg357_out;
SharedReg929_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg926_out;
   MUX_Product122_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg247_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg357_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg920_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg926_out_to_MUX_Product122_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_1_impl_0_out);

   Delay1No532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_1_impl_0_out,
                 Y => Delay1No532_out);

SharedReg918_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg933_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg933_out;
SharedReg852_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg852_out;
SharedReg851_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg851_out;
SharedReg814_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg814_out;
   MUX_Product122_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg933_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg852_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg851_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg814_out_to_MUX_Product122_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_1_impl_1_out);

   Delay1No533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_1_impl_1_out,
                 Y => Delay1No533_out);

Delay1No534_out_to_Product122_2_impl_parent_implementedSystem_port_0_cast <= Delay1No534_out;
Delay1No535_out_to_Product122_2_impl_parent_implementedSystem_port_1_cast <= Delay1No535_out;
   Product122_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_2_impl_out,
                 X => Delay1No534_out_to_Product122_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No535_out_to_Product122_2_impl_parent_implementedSystem_port_1_cast);

SharedReg926_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg926_out;
SharedReg93_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg93_out;
SharedReg250_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg250_out;
SharedReg520_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg520_out;
SharedReg929_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg920_out;
   MUX_Product122_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg926_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg250_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg520_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg920_out_to_MUX_Product122_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_2_impl_0_out);

   Delay1No534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_2_impl_0_out,
                 Y => Delay1No534_out);

SharedReg817_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg817_out;
SharedReg918_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg933_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg837_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg837_out;
SharedReg853_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg853_out;
   MUX_Product122_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg817_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg837_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg853_out_to_MUX_Product122_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_2_impl_1_out);

   Delay1No535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_2_impl_1_out,
                 Y => Delay1No535_out);

Delay1No536_out_to_Product122_3_impl_parent_implementedSystem_port_0_cast <= Delay1No536_out;
Delay1No537_out_to_Product122_3_impl_parent_implementedSystem_port_1_cast <= Delay1No537_out;
   Product122_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_3_impl_out,
                 X => Delay1No536_out_to_Product122_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No537_out_to_Product122_3_impl_parent_implementedSystem_port_1_cast);

SharedReg920_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg926_out;
SharedReg44_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg44_out;
SharedReg252_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg252_out;
SharedReg855_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg855_out;
SharedReg929_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product122_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg920_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg926_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg44_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg855_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product122_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_3_impl_0_out);

   Delay1No536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_3_impl_0_out,
                 Y => Delay1No536_out);

SharedReg855_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg855_out;
SharedReg820_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg820_out;
SharedReg918_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg933_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg933_out;
SharedReg821_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg821_out;
   MUX_Product122_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg855_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg820_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg933_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg821_out_to_MUX_Product122_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_3_impl_1_out);

   Delay1No537_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_3_impl_1_out,
                 Y => Delay1No537_out);

Delay1No538_out_to_Product122_4_impl_parent_implementedSystem_port_0_cast <= Delay1No538_out;
Delay1No539_out_to_Product122_4_impl_parent_implementedSystem_port_1_cast <= Delay1No539_out;
   Product122_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_4_impl_out,
                 X => Delay1No538_out_to_Product122_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No539_out_to_Product122_4_impl_parent_implementedSystem_port_1_cast);

SharedReg897_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg897_out;
SharedReg929_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg920_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg920_out;
SharedReg926_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg926_out;
SharedReg74_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg74_out;
SharedReg257_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg257_out;
   MUX_Product122_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg897_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg920_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg926_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg74_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg257_out_to_MUX_Product122_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_4_impl_0_out);

   Delay1No538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_4_impl_0_out,
                 Y => Delay1No538_out);

SharedReg933_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg933_out;
SharedReg857_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg857_out;
SharedReg898_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg898_out;
SharedReg843_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg843_out;
SharedReg918_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product122_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg933_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg857_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg898_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg843_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product122_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product122_4_impl_1_out);

   Delay1No539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_4_impl_1_out,
                 Y => Delay1No539_out);

Delay1No540_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast <= Delay1No540_out;
Delay1No541_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast <= Delay1No541_out;
   Product221_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_0_impl_out,
                 X => Delay1No540_out_to_Product221_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No541_out_to_Product221_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg908_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product221_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg922_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product221_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_0_impl_0_out);

   Delay1No540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_0_impl_0_out,
                 Y => Delay1No540_out);

SharedReg434_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg434_out;
SharedReg210_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg210_out;
SharedReg829_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg829_out;
SharedReg849_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg849_out;
SharedReg885_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg885_out;
SharedReg829_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg829_out;
   MUX_Product221_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg434_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg210_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg829_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg885_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg829_out_to_MUX_Product221_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_0_impl_1_out);

   Delay1No541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_0_impl_1_out,
                 Y => Delay1No541_out);

Delay1No542_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast <= Delay1No542_out;
Delay1No543_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast <= Delay1No543_out;
   Product221_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_1_impl_out,
                 X => Delay1No542_out_to_Product221_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No543_out_to_Product221_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg931_out;
   MUX_Product221_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg922_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg931_out_to_MUX_Product221_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_1_impl_0_out);

   Delay1No542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_1_impl_0_out,
                 Y => Delay1No542_out);

SharedReg833_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg833_out;
SharedReg438_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg438_out;
SharedReg214_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg214_out;
SharedReg833_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg833_out;
SharedReg832_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg832_out;
SharedReg887_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg887_out;
   MUX_Product221_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg833_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg438_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg214_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg833_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg832_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg887_out_to_MUX_Product221_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_1_impl_1_out);

   Delay1No543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_1_impl_1_out,
                 Y => Delay1No543_out);

Delay1No544_out_to_Product221_2_impl_parent_implementedSystem_port_0_cast <= Delay1No544_out;
Delay1No545_out_to_Product221_2_impl_parent_implementedSystem_port_1_cast <= Delay1No545_out;
   Product221_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_2_impl_out,
                 X => Delay1No544_out_to_Product221_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No545_out_to_Product221_2_impl_parent_implementedSystem_port_1_cast);

SharedReg931_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg931_out;
SharedReg908_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg922_out;
   MUX_Product221_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg931_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg922_out_to_MUX_Product221_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_2_impl_0_out);

   Delay1No544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_2_impl_0_out,
                 Y => Delay1No544_out);

SharedReg889_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg889_out;
SharedReg837_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg837_out;
SharedReg441_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg441_out;
SharedReg218_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg818_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg818_out;
SharedReg836_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg836_out;
   MUX_Product221_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg889_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg837_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg441_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg218_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg818_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg836_out_to_MUX_Product221_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_2_impl_1_out);

   Delay1No545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_2_impl_1_out,
                 Y => Delay1No545_out);

Delay1No546_out_to_Product221_3_impl_parent_implementedSystem_port_0_cast <= Delay1No546_out;
Delay1No547_out_to_Product221_3_impl_parent_implementedSystem_port_1_cast <= Delay1No547_out;
   Product221_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_3_impl_out,
                 X => Delay1No546_out_to_Product221_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No547_out_to_Product221_3_impl_parent_implementedSystem_port_1_cast);

SharedReg922_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg908_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product221_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg922_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product221_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_3_impl_0_out);

   Delay1No546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_3_impl_0_out,
                 Y => Delay1No546_out);

SharedReg840_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg840_out;
SharedReg891_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg891_out;
SharedReg841_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg841_out;
SharedReg411_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg222_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg222_out;
SharedReg892_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg892_out;
   MUX_Product221_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg840_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg891_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg841_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg222_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg892_out_to_MUX_Product221_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_3_impl_1_out);

   Delay1No547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_3_impl_1_out,
                 Y => Delay1No547_out);

Delay1No548_out_to_Product221_4_impl_parent_implementedSystem_port_0_cast <= Delay1No548_out;
Delay1No549_out_to_Product221_4_impl_parent_implementedSystem_port_1_cast <= Delay1No549_out;
   Product221_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_4_impl_out,
                 X => Delay1No548_out_to_Product221_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No549_out_to_Product221_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg908_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product221_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg922_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product221_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_4_impl_0_out);

   Delay1No548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_4_impl_0_out,
                 Y => Delay1No548_out);

SharedReg192_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg192_out;
SharedReg844_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg844_out;
SharedReg897_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg897_out;
SharedReg824_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg824_out;
SharedReg857_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg857_out;
SharedReg393_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg393_out;
   MUX_Product221_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg844_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg897_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg824_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg857_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg393_out_to_MUX_Product221_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product221_4_impl_1_out);

   Delay1No549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_4_impl_1_out,
                 Y => Delay1No549_out);

Delay1No550_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast <= Delay1No550_out;
Delay1No551_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast <= Delay1No551_out;
   Product321_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_0_impl_out,
                 X => Delay1No550_out_to_Product321_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No551_out_to_Product321_0_impl_parent_implementedSystem_port_1_cast);

SharedReg899_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg850_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg850_out;
SharedReg893_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg893_out;
SharedReg811_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg811_out;
SharedReg908_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product321_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg899_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg850_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg893_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg811_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product321_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_0_impl_0_out);

   Delay1No550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_0_out,
                 Y => Delay1No550_out);

SharedReg599_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg599_out;
SharedReg224_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg224_out;
SharedReg934_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg931_out;
SharedReg608_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg608_out;
   MUX_Product321_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg599_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg224_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg922_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg931_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg608_out_to_MUX_Product321_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_0_impl_1_out);

   Delay1No551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_0_impl_1_out,
                 Y => Delay1No551_out);

Delay1No552_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast <= Delay1No552_out;
Delay1No553_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast <= Delay1No553_out;
   Product321_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_1_impl_out,
                 X => Delay1No552_out_to_Product321_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No553_out_to_Product321_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg852_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg852_out;
SharedReg851_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg851_out;
SharedReg814_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg814_out;
   MUX_Product321_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg899_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg852_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg851_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg814_out_to_MUX_Product321_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_1_impl_0_out);

   Delay1No552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_0_out,
                 Y => Delay1No552_out);

SharedReg605_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg605_out;
SharedReg602_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg602_out;
SharedReg227_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg227_out;
SharedReg934_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg931_out;
   MUX_Product321_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg605_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg602_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg227_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg922_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg931_out_to_MUX_Product321_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_1_impl_1_out);

   Delay1No553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_1_impl_1_out,
                 Y => Delay1No553_out);

Delay1No554_out_to_Product321_2_impl_parent_implementedSystem_port_0_cast <= Delay1No554_out;
Delay1No555_out_to_Product321_2_impl_parent_implementedSystem_port_1_cast <= Delay1No555_out;
   Product321_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_2_impl_out,
                 X => Delay1No554_out_to_Product321_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No555_out_to_Product321_2_impl_parent_implementedSystem_port_1_cast);

SharedReg817_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg817_out;
SharedReg908_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg837_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg837_out;
SharedReg853_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg853_out;
   MUX_Product321_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg817_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg899_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg837_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg853_out_to_MUX_Product321_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_2_impl_0_out);

   Delay1No554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_2_impl_0_out,
                 Y => Delay1No554_out);

SharedReg931_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg931_out;
SharedReg444_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg444_out;
SharedReg614_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg614_out;
SharedReg232_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg934_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg922_out;
   MUX_Product321_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg931_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg444_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg614_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg922_out_to_MUX_Product321_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_2_impl_1_out);

   Delay1No555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_2_impl_1_out,
                 Y => Delay1No555_out);

Delay1No556_out_to_Product321_3_impl_parent_implementedSystem_port_0_cast <= Delay1No556_out;
Delay1No557_out_to_Product321_3_impl_parent_implementedSystem_port_1_cast <= Delay1No557_out;
   Product321_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_3_impl_out,
                 X => Delay1No556_out_to_Product321_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No557_out_to_Product321_3_impl_parent_implementedSystem_port_1_cast);

SharedReg855_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg855_out;
SharedReg820_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg820_out;
SharedReg908_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg899_out;
SharedReg900_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg821_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg821_out;
   MUX_Product321_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg855_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg820_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg899_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg821_out_to_MUX_Product321_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_3_impl_0_out);

   Delay1No556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_3_impl_0_out,
                 Y => Delay1No556_out);

SharedReg922_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg931_out;
SharedReg448_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg448_out;
SharedReg446_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg446_out;
SharedReg237_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg934_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product321_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg922_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg931_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg448_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg446_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product321_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_3_impl_1_out);

   Delay1No557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_3_impl_1_out,
                 Y => Delay1No557_out);

Delay1No558_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast <= Delay1No558_out;
Delay1No559_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast <= Delay1No559_out;
   Product321_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_4_impl_out,
                 X => Delay1No558_out_to_Product321_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No559_out_to_Product321_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg857_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg857_out;
SharedReg898_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg898_out;
SharedReg843_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg843_out;
SharedReg908_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg899_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg899_out;
   MUX_Product321_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg857_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg898_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg843_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg899_out_to_MUX_Product321_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_4_impl_0_out);

   Delay1No558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_4_impl_0_out,
                 Y => Delay1No558_out);

SharedReg242_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg242_out;
SharedReg934_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg922_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg922_out;
SharedReg931_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg931_out;
SharedReg634_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg634_out;
SharedReg450_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg450_out;
   MUX_Product321_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg242_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg922_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg931_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg634_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg450_out_to_MUX_Product321_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product321_4_impl_1_out);

   Delay1No559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_4_impl_1_out,
                 Y => Delay1No559_out);

Delay1No560_out_to_Subtract23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No560_out;
Delay1No561_out_to_Subtract23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No561_out;
   Subtract23_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract23_2_impl_out,
                 X => Delay1No560_out_to_Subtract23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No561_out_to_Subtract23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg262_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg262_out;
SharedReg643_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg643_out;
SharedReg14_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg611_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg611_out;
SharedReg149_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg149_out;
SharedReg342_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg342_out;
   MUX_Subtract23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg262_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg643_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg14_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg611_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg149_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg342_out_to_MUX_Subtract23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract23_2_impl_0_out);

   Delay1No560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_2_impl_0_out,
                 Y => Delay1No560_out);

SharedReg160_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg356_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg356_out;
SharedReg30_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg802_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg802_out;
SharedReg152_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg152_out;
SharedReg565_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg565_out;
   MUX_Subtract23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg356_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg30_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg802_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg565_out_to_MUX_Subtract23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract23_2_impl_1_out);

   Delay1No561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract23_2_impl_1_out,
                 Y => Delay1No561_out);

Delay1No562_out_to_Product124_0_impl_parent_implementedSystem_port_0_cast <= Delay1No562_out;
Delay1No563_out_to_Product124_0_impl_parent_implementedSystem_port_1_cast <= Delay1No563_out;
   Product124_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_0_impl_out,
                 X => Delay1No562_out_to_Product124_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No563_out_to_Product124_0_impl_parent_implementedSystem_port_1_cast);

SharedReg909_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg906_out;
SharedReg941_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg907_out;
SharedReg918_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product124_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg906_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg941_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg907_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product124_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_0_impl_0_out);

   Delay1No562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_0_impl_0_out,
                 Y => Delay1No562_out);

SharedReg434_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg434_out;
SharedReg210_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg210_out;
SharedReg33_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg33_out;
SharedReg636_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg636_out;
SharedReg108_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg108_out;
SharedReg829_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg829_out;
   MUX_Product124_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg434_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg210_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg33_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg636_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg108_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg829_out_to_MUX_Product124_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_0_impl_1_out);

   Delay1No563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_0_impl_1_out,
                 Y => Delay1No563_out);

Delay1No564_out_to_Product124_1_impl_parent_implementedSystem_port_0_cast <= Delay1No564_out;
Delay1No565_out_to_Product124_1_impl_parent_implementedSystem_port_1_cast <= Delay1No565_out;
   Product124_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_1_impl_out,
                 X => Delay1No564_out_to_Product124_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No565_out_to_Product124_1_impl_parent_implementedSystem_port_1_cast);

SharedReg918_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg906_out;
SharedReg941_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg907_out;
   MUX_Product124_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg906_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg941_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg907_out_to_MUX_Product124_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_1_impl_0_out);

   Delay1No564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_1_impl_0_out,
                 Y => Delay1No564_out);

SharedReg833_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg833_out;
SharedReg438_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg438_out;
SharedReg214_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg214_out;
SharedReg36_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
SharedReg624_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg624_out;
SharedReg124_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg124_out;
   MUX_Product124_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg833_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg438_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg214_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg624_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg124_out_to_MUX_Product124_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_1_impl_1_out);

   Delay1No565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_1_impl_1_out,
                 Y => Delay1No565_out);

Delay1No566_out_to_Product124_2_impl_parent_implementedSystem_port_0_cast <= Delay1No566_out;
Delay1No567_out_to_Product124_2_impl_parent_implementedSystem_port_1_cast <= Delay1No567_out;
   Product124_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_2_impl_out,
                 X => Delay1No566_out_to_Product124_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No567_out_to_Product124_2_impl_parent_implementedSystem_port_1_cast);

SharedReg907_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg907_out;
SharedReg918_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg941_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg941_out;
   MUX_Product124_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg907_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg941_out_to_MUX_Product124_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_2_impl_0_out);

   Delay1No566_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_2_impl_0_out,
                 Y => Delay1No566_out);

SharedReg113_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg113_out;
SharedReg837_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg837_out;
SharedReg441_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg441_out;
SharedReg218_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg218_out;
SharedReg91_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg91_out;
SharedReg645_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg645_out;
   MUX_Product124_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg837_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg441_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg218_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg91_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg645_out_to_MUX_Product124_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_2_impl_1_out);

   Delay1No567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_2_impl_1_out,
                 Y => Delay1No567_out);

Delay1No568_out_to_Product124_3_impl_parent_implementedSystem_port_0_cast <= Delay1No568_out;
Delay1No569_out_to_Product124_3_impl_parent_implementedSystem_port_1_cast <= Delay1No569_out;
   Product124_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_3_impl_out,
                 X => Delay1No568_out_to_Product124_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No569_out_to_Product124_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg907_out;
SharedReg918_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg906_out;
   MUX_Product124_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg907_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg906_out_to_MUX_Product124_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_3_impl_0_out);

   Delay1No568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_3_impl_0_out,
                 Y => Delay1No568_out);

SharedReg730_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg730_out;
SharedReg102_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg102_out;
SharedReg841_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg841_out;
SharedReg411_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg222_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg222_out;
SharedReg154_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg154_out;
   MUX_Product124_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg730_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg102_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg841_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg222_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_Product124_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_3_impl_1_out);

   Delay1No569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_3_impl_1_out,
                 Y => Delay1No569_out);

Delay1No570_out_to_Product124_4_impl_parent_implementedSystem_port_0_cast <= Delay1No570_out;
Delay1No571_out_to_Product124_4_impl_parent_implementedSystem_port_1_cast <= Delay1No571_out;
   Product124_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product124_4_impl_out,
                 X => Delay1No570_out_to_Product124_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No571_out_to_Product124_4_impl_parent_implementedSystem_port_1_cast);

SharedReg910_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg906_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg906_out;
SharedReg941_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg907_out;
SharedReg918_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product124_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg906_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg941_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg907_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product124_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_4_impl_0_out);

   Delay1No570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_4_impl_0_out,
                 Y => Delay1No570_out);

SharedReg192_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg192_out;
SharedReg46_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg46_out;
SharedReg754_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg754_out;
SharedReg98_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg98_out;
SharedReg857_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg857_out;
SharedReg393_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg393_out;
   MUX_Product124_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg46_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg754_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg98_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg857_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg393_out_to_MUX_Product124_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product124_4_impl_1_out);

   Delay1No571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product124_4_impl_1_out,
                 Y => Delay1No571_out);

Delay1No572_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast <= Delay1No572_out;
Delay1No573_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast <= Delay1No573_out;
   Product323_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_0_impl_out,
                 X => Delay1No572_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No573_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast);

SharedReg599_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg599_out;
SharedReg224_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg224_out;
SharedReg916_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg916_out;
SharedReg636_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg636_out;
SharedReg917_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg917_out;
SharedReg608_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg608_out;
   MUX_Product323_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg599_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg224_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg916_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg636_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg917_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg608_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_0_impl_0_out);

   Delay1No572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_0_impl_0_out,
                 Y => Delay1No572_out);

SharedReg909_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg33_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg33_out;
SharedReg945_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg945_out;
SharedReg108_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg108_out;
SharedReg918_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product323_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg909_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg33_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg108_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_0_impl_1_out);

   Delay1No573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_0_impl_1_out,
                 Y => Delay1No573_out);

Delay1No574_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast <= Delay1No574_out;
Delay1No575_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast <= Delay1No575_out;
   Product323_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_1_impl_out,
                 X => Delay1No574_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No575_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast);

SharedReg605_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg605_out;
SharedReg602_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg602_out;
SharedReg227_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg227_out;
SharedReg916_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg916_out;
SharedReg624_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg624_out;
SharedReg917_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg917_out;
   MUX_Product323_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg605_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg602_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg227_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg916_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg624_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg917_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_1_impl_0_out);

   Delay1No574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_1_impl_0_out,
                 Y => Delay1No574_out);

SharedReg918_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg36_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
SharedReg945_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg945_out;
SharedReg124_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg124_out;
   MUX_Product323_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg945_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg124_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_1_impl_1_out);

   Delay1No575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_1_impl_1_out,
                 Y => Delay1No575_out);

Delay1No576_out_to_Product323_2_impl_parent_implementedSystem_port_0_cast <= Delay1No576_out;
Delay1No577_out_to_Product323_2_impl_parent_implementedSystem_port_1_cast <= Delay1No577_out;
   Product323_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_2_impl_out,
                 X => Delay1No576_out_to_Product323_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No577_out_to_Product323_2_impl_parent_implementedSystem_port_1_cast);

SharedReg917_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg917_out;
SharedReg444_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg444_out;
SharedReg614_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg614_out;
SharedReg232_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg232_out;
SharedReg916_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg645_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg645_out;
   MUX_Product323_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg917_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg444_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg614_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg232_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg645_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_2_impl_0_out);

   Delay1No576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_2_impl_0_out,
                 Y => Delay1No576_out);

SharedReg113_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg113_out;
SharedReg918_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg91_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg91_out;
SharedReg945_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg945_out;
   MUX_Product323_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg113_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg909_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg91_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg945_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_2_impl_1_out);

   Delay1No577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_2_impl_1_out,
                 Y => Delay1No577_out);

Delay1No578_out_to_Product323_3_impl_parent_implementedSystem_port_0_cast <= Delay1No578_out;
Delay1No579_out_to_Product323_3_impl_parent_implementedSystem_port_1_cast <= Delay1No579_out;
   Product323_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_3_impl_out,
                 X => Delay1No578_out_to_Product323_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No579_out_to_Product323_3_impl_parent_implementedSystem_port_1_cast);

SharedReg730_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg730_out;
SharedReg917_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg917_out;
SharedReg448_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg448_out;
SharedReg446_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg446_out;
SharedReg237_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg916_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg916_out;
   MUX_Product323_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg730_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg917_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg448_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg446_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg916_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_3_impl_0_out);

   Delay1No578_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_3_impl_0_out,
                 Y => Delay1No578_out);

SharedReg945_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg945_out;
SharedReg102_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg102_out;
SharedReg918_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg909_out;
SharedReg910_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg154_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg154_out;
   MUX_Product323_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg945_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg102_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg909_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_3_impl_1_out);

   Delay1No579_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_3_impl_1_out,
                 Y => Delay1No579_out);

Delay1No580_out_to_Product323_4_impl_parent_implementedSystem_port_0_cast <= Delay1No580_out;
Delay1No581_out_to_Product323_4_impl_parent_implementedSystem_port_1_cast <= Delay1No581_out;
   Product323_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_4_impl_out,
                 X => Delay1No580_out_to_Product323_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No581_out_to_Product323_4_impl_parent_implementedSystem_port_1_cast);

SharedReg242_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg242_out;
SharedReg916_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg916_out;
SharedReg754_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg754_out;
SharedReg917_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg917_out;
SharedReg634_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg634_out;
SharedReg450_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg450_out;
   MUX_Product323_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg242_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg916_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg754_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg917_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg634_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg450_out_to_MUX_Product323_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_4_impl_0_out);

   Delay1No580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_4_impl_0_out,
                 Y => Delay1No580_out);

SharedReg910_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg46_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg46_out;
SharedReg945_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg945_out;
SharedReg98_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg98_out;
SharedReg918_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg909_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg909_out;
   MUX_Product323_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg46_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg945_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg98_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg909_out_to_MUX_Product323_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product323_4_impl_1_out);

   Delay1No581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_4_impl_1_out,
                 Y => Delay1No581_out);

Delay1No582_out_to_Subtract24_0_impl_parent_implementedSystem_port_0_cast <= Delay1No582_out;
Delay1No583_out_to_Subtract24_0_impl_parent_implementedSystem_port_1_cast <= Delay1No583_out;
   Subtract24_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_0_impl_out,
                 X => Delay1No582_out_to_Subtract24_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No583_out_to_Subtract24_0_impl_parent_implementedSystem_port_1_cast);

SharedReg663_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg663_out;
SharedReg5_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg570_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg570_out;
SharedReg210_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg210_out;
SharedReg600_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg600_out;
Delay3No215_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_6_cast <= Delay3No215_out;
   MUX_Subtract24_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg663_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg570_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg210_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg600_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No215_out_to_MUX_Subtract24_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_0_impl_0_out);

   Delay1No582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_0_impl_0_out,
                 Y => Delay1No582_out);

SharedReg688_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg688_out;
SharedReg21_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg707_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg707_out;
SharedReg211_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg211_out;
SharedReg402_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg402_out;
Delay3No220_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_6_cast <= Delay3No220_out;
   MUX_Subtract24_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg688_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg707_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg211_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg402_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No220_out_to_MUX_Subtract24_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_0_impl_1_out);

   Delay1No583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_0_impl_1_out,
                 Y => Delay1No583_out);

Delay1No584_out_to_Subtract24_1_impl_parent_implementedSystem_port_0_cast <= Delay1No584_out;
Delay1No585_out_to_Subtract24_1_impl_parent_implementedSystem_port_1_cast <= Delay1No585_out;
   Subtract24_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_1_impl_out,
                 X => Delay1No584_out_to_Subtract24_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No585_out_to_Subtract24_1_impl_parent_implementedSystem_port_1_cast);

Delay3No216_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No216_out;
SharedReg665_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg665_out;
SharedReg5_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg573_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg573_out;
SharedReg604_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg604_out;
SharedReg279_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg279_out;
   MUX_Subtract24_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No216_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg665_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg573_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg604_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg279_out_to_MUX_Subtract24_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_1_impl_0_out);

   Delay1No584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_1_impl_0_out,
                 Y => Delay1No584_out);

Delay3No221_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_1_cast <= Delay3No221_out;
SharedReg689_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg689_out;
SharedReg21_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg709_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg709_out;
SharedReg744_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg744_out;
SharedReg213_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg213_out;
   MUX_Subtract24_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No221_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg689_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg21_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg709_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg744_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg213_out_to_MUX_Subtract24_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_1_impl_1_out);

   Delay1No585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_1_impl_1_out,
                 Y => Delay1No585_out);

Delay1No586_out_to_Subtract24_2_impl_parent_implementedSystem_port_0_cast <= Delay1No586_out;
Delay1No587_out_to_Subtract24_2_impl_parent_implementedSystem_port_1_cast <= Delay1No587_out;
   Subtract24_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_2_impl_out,
                 X => Delay1No586_out_to_Subtract24_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No587_out_to_Subtract24_2_impl_parent_implementedSystem_port_1_cast);

SharedReg442_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg442_out;
SharedReg504_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg504_out;
SharedReg554_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg554_out;
SharedReg4_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg4_out;
SharedReg576_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg576_out;
SharedReg443_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg443_out;
   MUX_Subtract24_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg442_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg504_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg554_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg576_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg443_out_to_MUX_Subtract24_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_2_impl_0_out);

   Delay1No586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_2_impl_0_out,
                 Y => Delay1No586_out);

SharedReg408_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg408_out;
SharedReg564_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg564_out;
SharedReg589_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg589_out;
SharedReg20_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg20_out;
SharedReg711_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg711_out;
SharedReg747_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg747_out;
   MUX_Subtract24_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg408_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg564_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg589_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg20_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg711_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg747_out_to_MUX_Subtract24_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_2_impl_1_out);

   Delay1No587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_2_impl_1_out,
                 Y => Delay1No587_out);

Delay1No588_out_to_Subtract24_3_impl_parent_implementedSystem_port_0_cast <= Delay1No588_out;
Delay1No589_out_to_Subtract24_3_impl_parent_implementedSystem_port_1_cast <= Delay1No589_out;
   Subtract24_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_3_impl_out,
                 X => Delay1No588_out_to_Subtract24_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No589_out_to_Subtract24_3_impl_parent_implementedSystem_port_1_cast);

SharedReg206_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg206_out;
SharedReg268_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg268_out;
Delay3No198_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_3_cast <= Delay3No198_out;
SharedReg486_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg486_out;
SharedReg4_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg579_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg579_out;
   MUX_Subtract24_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg206_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg268_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No198_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg486_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg4_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg579_out_to_MUX_Subtract24_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_3_impl_0_out);

   Delay1No588_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_3_impl_0_out,
                 Y => Delay1No588_out);

SharedReg207_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg45_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg45_out;
Delay3No213_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_3_cast <= Delay3No213_out;
SharedReg516_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg516_out;
SharedReg20_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg713_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg713_out;
   MUX_Subtract24_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg45_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No213_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg516_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg713_out_to_MUX_Subtract24_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_3_impl_1_out);

   Delay1No589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_3_impl_1_out,
                 Y => Delay1No589_out);

Delay1No590_out_to_Subtract24_4_impl_parent_implementedSystem_port_0_cast <= Delay1No590_out;
Delay1No591_out_to_Subtract24_4_impl_parent_implementedSystem_port_1_cast <= Delay1No591_out;
   Subtract24_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_4_impl_out,
                 X => Delay1No590_out_to_Subtract24_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No591_out_to_Subtract24_4_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg582_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg582_out;
SharedReg399_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg399_out;
SharedReg632_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg632_out;
SharedReg508_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg508_out;
SharedReg671_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg671_out;
   MUX_Subtract24_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg582_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg399_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg632_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg508_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg671_out_to_MUX_Subtract24_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_4_impl_0_out);

   Delay1No590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_4_impl_0_out,
                 Y => Delay1No590_out);

SharedReg21_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg715_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg715_out;
SharedReg334_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg334_out;
SharedReg862_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg862_out;
SharedReg568_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg568_out;
SharedReg692_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg692_out;
   MUX_Subtract24_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg715_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg334_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg862_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg568_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg692_out_to_MUX_Subtract24_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract24_4_impl_1_out);

   Delay1No591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_4_impl_1_out,
                 Y => Delay1No591_out);

Delay1No592_out_to_Subtract26_0_impl_parent_implementedSystem_port_0_cast <= Delay1No592_out;
Delay1No593_out_to_Subtract26_0_impl_parent_implementedSystem_port_1_cast <= Delay1No593_out;
   Subtract26_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_0_impl_out,
                 X => Delay1No592_out_to_Subtract26_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No593_out_to_Subtract26_0_impl_parent_implementedSystem_port_1_cast);

SharedReg245_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg245_out;
SharedReg6_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg663_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg663_out;
SharedReg601_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg601_out;
SharedReg523_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg523_out;
SharedReg683_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg683_out;
   MUX_Subtract26_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg245_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg663_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg601_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg523_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg683_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_0_impl_0_out);

   Delay1No592_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_0_impl_0_out,
                 Y => Delay1No592_out);

SharedReg261_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg22_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg688_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg688_out;
SharedReg740_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg740_out;
SharedReg209_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg209_out;
SharedReg706_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg706_out;
   MUX_Subtract26_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg688_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg740_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg209_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg706_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_0_impl_1_out);

   Delay1No593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_0_impl_1_out,
                 Y => Delay1No593_out);

Delay1No594_out_to_Subtract26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No594_out;
Delay1No595_out_to_Subtract26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No595_out;
   Subtract26_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_1_impl_out,
                 X => Delay1No594_out_to_Subtract26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No595_out_to_Subtract26_1_impl_parent_implementedSystem_port_1_cast);

SharedReg684_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg684_out;
SharedReg248_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg248_out;
SharedReg6_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg665_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg665_out;
SharedReg249_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg249_out;
SharedReg603_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg603_out;
   MUX_Subtract26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg684_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg248_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg6_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg665_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg249_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg603_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_1_impl_0_out);

   Delay1No594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_1_impl_0_out,
                 Y => Delay1No594_out);

SharedReg708_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg708_out;
SharedReg264_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg22_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg689_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg689_out;
SharedReg150_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg150_out;
SharedReg438_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg438_out;
   MUX_Subtract26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg708_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg22_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg689_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg150_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg438_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_1_impl_1_out);

   Delay1No595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_1_impl_1_out,
                 Y => Delay1No595_out);

Delay1No596_out_to_Subtract26_2_impl_parent_implementedSystem_port_0_cast <= Delay1No596_out;
Delay1No597_out_to_Subtract26_2_impl_parent_implementedSystem_port_1_cast <= Delay1No597_out;
   Subtract26_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_2_impl_out,
                 X => Delay1No596_out_to_Subtract26_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No597_out_to_Subtract26_2_impl_parent_implementedSystem_port_1_cast);

SharedReg282_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg282_out;
Delay3No217_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_2_cast <= Delay3No217_out;
SharedReg667_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg667_out;
SharedReg5_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg5_out;
SharedReg667_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg667_out;
SharedReg233_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg233_out;
   MUX_Subtract26_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No217_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg667_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg5_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg667_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg233_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_2_impl_0_out);

   Delay1No596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_2_impl_0_out,
                 Y => Delay1No596_out);

SharedReg217_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg217_out;
Delay3No222_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_2_cast <= Delay3No222_out;
SharedReg690_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg690_out;
SharedReg21_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
SharedReg690_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg690_out;
SharedReg532_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg532_out;
   MUX_Subtract26_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg217_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No222_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg690_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg690_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg532_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_2_impl_1_out);

   Delay1No597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_2_impl_1_out,
                 Y => Delay1No597_out);

Delay1No598_out_to_Subtract26_3_impl_parent_implementedSystem_port_0_cast <= Delay1No598_out;
Delay1No599_out_to_Subtract26_3_impl_parent_implementedSystem_port_1_cast <= Delay1No599_out;
   Subtract26_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_3_impl_out,
                 X => Delay1No598_out_to_Subtract26_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No599_out_to_Subtract26_3_impl_parent_implementedSystem_port_1_cast);

SharedReg413_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg413_out;
SharedReg447_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg447_out;
SharedReg506_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg506_out;
SharedReg556_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg556_out;
SharedReg5_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg669_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg669_out;
   MUX_Subtract26_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg413_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg447_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg506_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg556_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg669_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_3_impl_0_out);

   Delay1No598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_3_impl_0_out,
                 Y => Delay1No598_out);

SharedReg751_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg751_out;
SharedReg411_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg411_out;
SharedReg566_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg591_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg591_out;
SharedReg21_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg691_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg691_out;
   MUX_Subtract26_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg751_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg411_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg566_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg591_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg691_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_3_impl_1_out);

   Delay1No599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_3_impl_1_out,
                 Y => Delay1No599_out);

Delay1No600_out_to_Subtract26_4_impl_parent_implementedSystem_port_0_cast <= Delay1No600_out;
Delay1No601_out_to_Subtract26_4_impl_parent_implementedSystem_port_1_cast <= Delay1No601_out;
   Subtract26_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_4_impl_out,
                 X => Delay1No600_out_to_Subtract26_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No601_out_to_Subtract26_4_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg671_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg671_out;
SharedReg242_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg242_out;
SharedReg270_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg270_out;
Delay3No219_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_5_cast <= Delay3No219_out;
SharedReg258_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg258_out;
   MUX_Subtract26_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg671_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg242_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg270_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No219_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg258_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_4_impl_0_out);

   Delay1No600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_4_impl_0_out,
                 Y => Delay1No600_out);

SharedReg22_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg692_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg692_out;
SharedReg193_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg193_out;
SharedReg660_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg660_out;
Delay3No224_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_5_cast <= Delay3No224_out;
SharedReg273_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg273_out;
   MUX_Subtract26_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg692_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg193_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg660_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay3No224_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg273_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract26_4_impl_1_out);

   Delay1No601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_4_impl_1_out,
                 Y => Delay1No601_out);

Delay1No602_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast <= Delay1No602_out;
Delay1No603_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast <= Delay1No603_out;
   Product55_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_0_impl_out,
                 X => Delay1No602_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No603_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast);

SharedReg949_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg929_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg929_out;
SharedReg941_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product55_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg949_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg929_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg941_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg907_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_0_impl_0_out);

   Delay1No602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_0_impl_0_out,
                 Y => Delay1No602_out);

SharedReg606_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg606_out;
SharedReg259_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg259_out;
SharedReg894_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg894_out;
SharedReg875_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg875_out;
SharedReg637_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg637_out;
SharedReg719_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg719_out;
   MUX_Product55_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg606_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg259_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg894_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg875_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg637_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg719_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_0_impl_1_out);

   Delay1No603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_0_impl_1_out,
                 Y => Delay1No603_out);

Delay1No604_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast <= Delay1No604_out;
Delay1No605_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast <= Delay1No605_out;
   Product55_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_1_impl_out,
                 X => Delay1No604_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No605_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg949_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg929_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg929_out;
SharedReg941_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg907_out;
   MUX_Product55_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg949_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg929_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg941_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg907_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_1_impl_0_out);

   Delay1No604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_1_impl_0_out,
                 Y => Delay1No604_out);

SharedReg642_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg642_out;
SharedReg610_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg610_out;
SharedReg262_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg262_out;
SharedReg694_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg694_out;
SharedReg867_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg867_out;
SharedReg626_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg626_out;
   MUX_Product55_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg642_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg610_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg262_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg694_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg867_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg626_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_1_impl_1_out);

   Delay1No605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_1_impl_1_out,
                 Y => Delay1No605_out);

Delay1No606_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast <= Delay1No606_out;
Delay1No607_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast <= Delay1No607_out;
   Product55_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_2_impl_out,
                 X => Delay1No606_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No607_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast);

SharedReg907_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg949_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg929_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg941_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg941_out;
   MUX_Product55_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg907_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg949_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg941_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_2_impl_0_out);

   Delay1No606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_2_impl_0_out,
                 Y => Delay1No606_out);

SharedReg630_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg630_out;
SharedReg647_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg647_out;
SharedReg628_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg628_out;
SharedReg265_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg265_out;
SharedReg854_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg854_out;
SharedReg869_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg869_out;
   MUX_Product55_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg630_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg647_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg628_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg265_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg854_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg869_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_2_impl_1_out);

   Delay1No607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_2_impl_1_out,
                 Y => Delay1No607_out);

Delay1No608_out_to_Product55_3_impl_parent_implementedSystem_port_0_cast <= Delay1No608_out;
Delay1No609_out_to_Product55_3_impl_parent_implementedSystem_port_1_cast <= Delay1No609_out;
   Product55_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_3_impl_out,
                 X => Delay1No608_out_to_Product55_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No609_out_to_Product55_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg949_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg929_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg929_out;
   MUX_Product55_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg907_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg949_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg929_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_3_impl_0_out);

   Delay1No608_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_3_impl_0_out,
                 Y => Delay1No608_out);

SharedReg871_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg871_out;
SharedReg652_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg652_out;
SharedReg732_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg732_out;
SharedReg617_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg617_out;
SharedReg269_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg269_out;
SharedReg841_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg841_out;
   MUX_Product55_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg871_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg652_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg732_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg617_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg269_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg841_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_3_impl_1_out);

   Delay1No609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_3_impl_1_out,
                 Y => Delay1No609_out);

Delay1No610_out_to_Product55_4_impl_parent_implementedSystem_port_0_cast <= Delay1No610_out;
Delay1No611_out_to_Product55_4_impl_parent_implementedSystem_port_1_cast <= Delay1No611_out;
   Product55_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_4_impl_out,
                 X => Delay1No610_out_to_Product55_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No611_out_to_Product55_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg929_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg929_out;
SharedReg941_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg941_out;
SharedReg907_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg949_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg949_out;
   MUX_Product55_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg929_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg941_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg907_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg949_out_to_MUX_Product55_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_4_impl_0_out);

   Delay1No610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_4_impl_0_out,
                 Y => Delay1No610_out);

SharedReg271_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg896_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg896_out;
SharedReg824_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg824_out;
SharedReg736_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg736_out;
SharedReg757_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg757_out;
SharedReg595_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
   MUX_Product55_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg896_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg824_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg736_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg757_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Product55_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product55_4_impl_1_out);

   Delay1No611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_4_impl_1_out,
                 Y => Delay1No611_out);

Delay1No612_out_to_Product127_0_impl_parent_implementedSystem_port_0_cast <= Delay1No612_out;
Delay1No613_out_to_Product127_0_impl_parent_implementedSystem_port_1_cast <= Delay1No613_out;
   Product127_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_0_impl_out,
                 X => Delay1No612_out_to_Product127_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No613_out_to_Product127_0_impl_parent_implementedSystem_port_1_cast);

SharedReg949_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg934_out;
SharedReg941_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg941_out;
SharedReg917_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg917_out;
SharedReg719_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg719_out;
   MUX_Product127_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg949_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg900_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg934_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg941_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg917_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg719_out_to_MUX_Product127_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_0_impl_0_out);

   Delay1No612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_0_impl_0_out,
                 Y => Delay1No612_out);

SharedReg620_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg620_out;
SharedReg275_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg894_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg894_out;
SharedReg885_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg885_out;
SharedReg637_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg637_out;
SharedReg918_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product127_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg620_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg894_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg885_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg637_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product127_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_0_impl_1_out);

   Delay1No613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_0_impl_1_out,
                 Y => Delay1No613_out);

Delay1No614_out_to_Product127_1_impl_parent_implementedSystem_port_0_cast <= Delay1No614_out;
Delay1No615_out_to_Product127_1_impl_parent_implementedSystem_port_1_cast <= Delay1No615_out;
   Product127_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_1_impl_out,
                 X => Delay1No614_out_to_Product127_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No615_out_to_Product127_1_impl_parent_implementedSystem_port_1_cast);

SharedReg642_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg642_out;
SharedReg949_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg934_out;
SharedReg941_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg941_out;
SharedReg917_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg917_out;
   MUX_Product127_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg642_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg949_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg934_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg941_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg917_out_to_MUX_Product127_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_1_impl_0_out);

   Delay1No614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_1_impl_0_out,
                 Y => Delay1No614_out);

SharedReg918_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg624_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg624_out;
SharedReg279_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg279_out;
SharedReg694_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg694_out;
SharedReg877_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg877_out;
SharedReg626_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg626_out;
   MUX_Product127_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg624_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg279_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg694_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg877_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg626_out_to_MUX_Product127_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_1_impl_1_out);

   Delay1No615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_1_impl_1_out,
                 Y => Delay1No615_out);

Delay1No616_out_to_Product127_2_impl_parent_implementedSystem_port_0_cast <= Delay1No616_out;
Delay1No617_out_to_Product127_2_impl_parent_implementedSystem_port_1_cast <= Delay1No617_out;
   Product127_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_2_impl_out,
                 X => Delay1No616_out_to_Product127_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No617_out_to_Product127_2_impl_parent_implementedSystem_port_1_cast);

SharedReg917_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg917_out;
SharedReg647_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg647_out;
SharedReg949_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg934_out;
SharedReg941_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg941_out;
   MUX_Product127_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg917_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg647_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg949_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg900_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg934_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg941_out_to_MUX_Product127_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_2_impl_0_out);

   Delay1No616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_2_impl_0_out,
                 Y => Delay1No616_out);

SharedReg630_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg630_out;
SharedReg918_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg645_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg645_out;
SharedReg282_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg282_out;
SharedReg854_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg854_out;
SharedReg879_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg879_out;
   MUX_Product127_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg630_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg645_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg282_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg854_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg879_out_to_MUX_Product127_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_2_impl_1_out);

   Delay1No617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_2_impl_1_out,
                 Y => Delay1No617_out);

Delay1No618_out_to_Product127_3_impl_parent_implementedSystem_port_0_cast <= Delay1No618_out;
Delay1No619_out_to_Product127_3_impl_parent_implementedSystem_port_1_cast <= Delay1No619_out;
   Product127_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_3_impl_out,
                 X => Delay1No618_out_to_Product127_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No619_out_to_Product127_3_impl_parent_implementedSystem_port_1_cast);

SharedReg941_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg941_out;
SharedReg917_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg917_out;
SharedReg732_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg732_out;
SharedReg949_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg949_out;
SharedReg900_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg934_out;
   MUX_Product127_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg941_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg917_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg732_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg949_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg900_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg934_out_to_MUX_Product127_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_3_impl_0_out);

   Delay1No618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_3_impl_0_out,
                 Y => Delay1No618_out);

SharedReg881_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg881_out;
SharedReg652_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg652_out;
SharedReg918_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg650_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg650_out;
SharedReg284_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg841_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg841_out;
   MUX_Product127_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg881_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg652_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg650_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg841_out_to_MUX_Product127_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_3_impl_1_out);

   Delay1No619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_3_impl_1_out,
                 Y => Delay1No619_out);

Delay1No620_out_to_Product127_4_impl_parent_implementedSystem_port_0_cast <= Delay1No620_out;
Delay1No621_out_to_Product127_4_impl_parent_implementedSystem_port_1_cast <= Delay1No621_out;
   Product127_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_4_impl_out,
                 X => Delay1No620_out_to_Product127_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No621_out_to_Product127_4_impl_parent_implementedSystem_port_1_cast);

SharedReg900_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg900_out;
SharedReg934_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg934_out;
SharedReg941_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg941_out;
SharedReg917_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg917_out;
SharedReg757_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg757_out;
SharedReg949_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg949_out;
   MUX_Product127_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg900_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg934_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg941_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg917_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg757_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg949_out_to_MUX_Product127_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_4_impl_0_out);

   Delay1No620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_4_impl_0_out,
                 Y => Delay1No620_out);

SharedReg287_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg287_out;
SharedReg896_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg896_out;
SharedReg843_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg843_out;
SharedReg736_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg736_out;
SharedReg918_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg632_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg632_out;
   MUX_Product127_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg287_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg896_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg843_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg736_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg632_out_to_MUX_Product127_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product127_4_impl_1_out);

   Delay1No621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_4_impl_1_out,
                 Y => Delay1No621_out);

Delay1No622_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast <= Delay1No622_out;
Delay1No623_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast <= Delay1No623_out;
   Product226_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_0_impl_out,
                 X => Delay1No622_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No623_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast);

SharedReg950_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg901_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg901_out;
SharedReg945_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg945_out;
SharedReg907_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg908_out;
   MUX_Product226_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg950_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg901_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg907_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg908_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_0_impl_0_out);

   Delay1No622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_0_impl_0_out,
                 Y => Delay1No622_out);

SharedReg606_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg606_out;
SharedReg259_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg259_out;
SharedReg121_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg121_out;
SharedReg875_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg875_out;
SharedReg800_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg741_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg741_out;
   MUX_Product226_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg606_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg259_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg121_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg875_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg741_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_0_impl_1_out);

   Delay1No623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_0_impl_1_out,
                 Y => Delay1No623_out);

Delay1No624_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast <= Delay1No624_out;
Delay1No625_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast <= Delay1No625_out;
   Product226_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_1_impl_out,
                 X => Delay1No624_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No625_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast);

SharedReg908_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg908_out;
SharedReg950_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg901_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg901_out;
SharedReg945_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg945_out;
SharedReg907_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg907_out;
   MUX_Product226_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg908_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg950_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg901_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg945_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg907_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_1_impl_0_out);

   Delay1No624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_1_impl_0_out,
                 Y => Delay1No624_out);

SharedReg724_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg724_out;
SharedReg610_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg610_out;
SharedReg262_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg262_out;
SharedReg138_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg138_out;
SharedReg867_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg867_out;
SharedReg744_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg744_out;
   MUX_Product226_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg724_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg610_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg262_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg138_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg867_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg744_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_1_impl_1_out);

   Delay1No625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_1_impl_1_out,
                 Y => Delay1No625_out);

Delay1No626_out_to_Product226_2_impl_parent_implementedSystem_port_0_cast <= Delay1No626_out;
Delay1No627_out_to_Product226_2_impl_parent_implementedSystem_port_1_cast <= Delay1No627_out;
   Product226_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_2_impl_out,
                 X => Delay1No626_out_to_Product226_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No627_out_to_Product226_2_impl_parent_implementedSystem_port_1_cast);

SharedReg907_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg908_out;
SharedReg950_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg901_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg901_out;
SharedReg945_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg945_out;
   MUX_Product226_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg907_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg908_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg950_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg901_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg945_out_to_MUX_Product226_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_2_impl_0_out);

   Delay1No626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_2_impl_0_out,
                 Y => Delay1No626_out);

SharedReg747_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg747_out;
SharedReg728_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg728_out;
SharedReg628_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg628_out;
SharedReg265_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg265_out;
SharedReg141_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg141_out;
SharedReg869_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg869_out;
   MUX_Product226_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg747_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg728_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg628_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg265_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg141_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg869_out_to_MUX_Product226_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_2_impl_1_out);

   Delay1No627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_2_impl_1_out,
                 Y => Delay1No627_out);

Delay1No628_out_to_Product226_3_impl_parent_implementedSystem_port_0_cast <= Delay1No628_out;
Delay1No629_out_to_Product226_3_impl_parent_implementedSystem_port_1_cast <= Delay1No629_out;
   Product226_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_3_impl_out,
                 X => Delay1No628_out_to_Product226_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No629_out_to_Product226_3_impl_parent_implementedSystem_port_1_cast);

SharedReg945_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg945_out;
SharedReg907_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg908_out;
SharedReg950_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg901_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg901_out;
   MUX_Product226_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg945_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg907_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg908_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg950_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg901_out_to_MUX_Product226_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_3_impl_0_out);

   Delay1No628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_3_impl_0_out,
                 Y => Delay1No628_out);

SharedReg871_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg871_out;
SharedReg806_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg806_out;
SharedReg752_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg617_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg617_out;
SharedReg269_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg269_out;
SharedReg129_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg129_out;
   MUX_Product226_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg871_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg806_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg617_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg269_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg129_out_to_MUX_Product226_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_3_impl_1_out);

   Delay1No629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_3_impl_1_out,
                 Y => Delay1No629_out);

Delay1No630_out_to_Product226_4_impl_parent_implementedSystem_port_0_cast <= Delay1No630_out;
Delay1No631_out_to_Product226_4_impl_parent_implementedSystem_port_1_cast <= Delay1No631_out;
   Product226_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_4_impl_out,
                 X => Delay1No630_out_to_Product226_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No631_out_to_Product226_4_impl_parent_implementedSystem_port_1_cast);

SharedReg910_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg901_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg901_out;
SharedReg945_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg945_out;
SharedReg907_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg907_out;
SharedReg908_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg908_out;
SharedReg950_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg950_out;
   MUX_Product226_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg901_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg945_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg907_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg908_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg950_out_to_MUX_Product226_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_4_impl_0_out);

   Delay1No630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_4_impl_0_out,
                 Y => Delay1No630_out);

SharedReg271_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg105_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg824_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg824_out;
SharedReg864_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg864_out;
SharedReg810_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg810_out;
SharedReg595_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
   MUX_Product226_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg824_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg864_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg810_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Product226_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product226_4_impl_1_out);

   Delay1No631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_4_impl_1_out,
                 Y => Delay1No631_out);

Delay1No632_out_to_Product326_0_impl_parent_implementedSystem_port_0_cast <= Delay1No632_out;
Delay1No633_out_to_Product326_0_impl_parent_implementedSystem_port_1_cast <= Delay1No633_out;
   Product326_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_0_impl_out,
                 X => Delay1No632_out_to_Product326_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No633_out_to_Product326_0_impl_parent_implementedSystem_port_1_cast);

SharedReg620_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg620_out;
SharedReg275_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg911_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg911_out;
SharedReg885_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg885_out;
SharedReg800_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg918_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
   MUX_Product326_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg620_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg911_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg885_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Product326_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_0_impl_0_out);

   Delay1No632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_0_impl_0_out,
                 Y => Delay1No632_out);

SharedReg950_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg121_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg121_out;
SharedReg945_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg945_out;
SharedReg917_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg917_out;
SharedReg741_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg741_out;
   MUX_Product326_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg950_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg121_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg945_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg917_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg741_out_to_MUX_Product326_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_0_impl_1_out);

   Delay1No633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_0_impl_1_out,
                 Y => Delay1No633_out);

Delay1No634_out_to_Product326_1_impl_parent_implementedSystem_port_0_cast <= Delay1No634_out;
Delay1No635_out_to_Product326_1_impl_parent_implementedSystem_port_1_cast <= Delay1No635_out;
   Product326_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_1_impl_out,
                 X => Delay1No634_out_to_Product326_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No635_out_to_Product326_1_impl_parent_implementedSystem_port_1_cast);

SharedReg918_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg918_out;
SharedReg624_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg624_out;
SharedReg279_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg279_out;
SharedReg911_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg911_out;
SharedReg877_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg877_out;
SharedReg744_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg744_out;
   MUX_Product326_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg918_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg624_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg279_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg911_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg877_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg744_out_to_MUX_Product326_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_1_impl_0_out);

   Delay1No634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_1_impl_0_out,
                 Y => Delay1No634_out);

SharedReg724_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg724_out;
SharedReg950_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg910_out;
SharedReg138_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg138_out;
SharedReg945_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg945_out;
SharedReg917_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg917_out;
   MUX_Product326_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg724_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg950_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg910_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg138_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg945_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg917_out_to_MUX_Product326_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_1_impl_1_out);

   Delay1No635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_1_impl_1_out,
                 Y => Delay1No635_out);

Delay1No636_out_to_Product326_2_impl_parent_implementedSystem_port_0_cast <= Delay1No636_out;
Delay1No637_out_to_Product326_2_impl_parent_implementedSystem_port_1_cast <= Delay1No637_out;
   Product326_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_2_impl_out,
                 X => Delay1No636_out_to_Product326_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No637_out_to_Product326_2_impl_parent_implementedSystem_port_1_cast);

SharedReg747_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg747_out;
SharedReg918_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg918_out;
SharedReg645_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg645_out;
SharedReg282_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg282_out;
SharedReg911_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg911_out;
SharedReg879_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg879_out;
   MUX_Product326_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg747_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg918_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg645_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg282_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg911_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg879_out_to_MUX_Product326_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_2_impl_0_out);

   Delay1No636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_2_impl_0_out,
                 Y => Delay1No636_out);

SharedReg917_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg917_out;
SharedReg728_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg728_out;
SharedReg950_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg910_out;
SharedReg141_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg141_out;
SharedReg945_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg945_out;
   MUX_Product326_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg917_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg728_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg950_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg910_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg141_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg945_out_to_MUX_Product326_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_2_impl_1_out);

   Delay1No637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_2_impl_1_out,
                 Y => Delay1No637_out);

Delay1No638_out_to_Product326_3_impl_parent_implementedSystem_port_0_cast <= Delay1No638_out;
Delay1No639_out_to_Product326_3_impl_parent_implementedSystem_port_1_cast <= Delay1No639_out;
   Product326_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_3_impl_out,
                 X => Delay1No638_out_to_Product326_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No639_out_to_Product326_3_impl_parent_implementedSystem_port_1_cast);

SharedReg881_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg881_out;
SharedReg806_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg806_out;
SharedReg918_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg918_out;
SharedReg650_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg650_out;
SharedReg284_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg911_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg911_out;
   MUX_Product326_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg881_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg806_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg918_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg650_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg911_out_to_MUX_Product326_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_3_impl_0_out);

   Delay1No638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_3_impl_0_out,
                 Y => Delay1No638_out);

SharedReg945_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg945_out;
SharedReg917_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg917_out;
SharedReg752_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg950_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg950_out;
SharedReg910_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg910_out;
SharedReg129_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg129_out;
   MUX_Product326_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg945_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg917_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg950_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg910_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg129_out_to_MUX_Product326_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_3_impl_1_out);

   Delay1No639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_3_impl_1_out,
                 Y => Delay1No639_out);

Delay1No640_out_to_Product326_4_impl_parent_implementedSystem_port_0_cast <= Delay1No640_out;
Delay1No641_out_to_Product326_4_impl_parent_implementedSystem_port_1_cast <= Delay1No641_out;
   Product326_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_4_impl_out,
                 X => Delay1No640_out_to_Product326_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No641_out_to_Product326_4_impl_parent_implementedSystem_port_1_cast);

SharedReg287_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg287_out;
SharedReg911_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg911_out;
SharedReg843_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg843_out;
SharedReg864_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg864_out;
SharedReg918_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg918_out;
SharedReg632_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg632_out;
   MUX_Product326_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg287_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg911_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg843_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg864_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg918_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg632_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_4_impl_0_out);

   Delay1No640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_4_impl_0_out,
                 Y => Delay1No640_out);

SharedReg910_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg910_out;
SharedReg105_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg945_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg945_out;
SharedReg917_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg917_out;
SharedReg810_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg810_out;
SharedReg950_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg950_out;
   MUX_Product326_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg910_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg945_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg917_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg810_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg950_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Product326_4_impl_1_out);

   Delay1No641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_4_impl_1_out,
                 Y => Delay1No641_out);

Delay1No642_out_to_Subtract27_0_impl_parent_implementedSystem_port_0_cast <= Delay1No642_out;
Delay1No643_out_to_Subtract27_0_impl_parent_implementedSystem_port_1_cast <= Delay1No643_out;
   Subtract27_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract27_0_impl_out,
                 X => Delay1No642_out_to_Subtract27_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No643_out_to_Subtract27_0_impl_parent_implementedSystem_port_1_cast);

SharedReg403_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg403_out;
SharedReg7_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg759_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg759_out;
SharedReg246_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg246_out;
SharedReg607_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg607_out;
SharedReg758_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg758_out;
   MUX_Subtract27_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg403_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg759_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg246_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg607_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg758_out_to_MUX_Subtract27_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_0_impl_0_out);

   Delay1No642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_0_impl_0_out,
                 Y => Delay1No642_out);

SharedReg437_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg437_out;
SharedReg23_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg789_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg789_out;
SharedReg540_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg540_out;
SharedReg434_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg434_out;
SharedReg788_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg788_out;
   MUX_Subtract27_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg437_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg789_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg540_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg434_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg788_out_to_MUX_Subtract27_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_0_impl_1_out);

   Delay1No643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_0_impl_1_out,
                 Y => Delay1No643_out);

Delay1No644_out_to_Subtract27_1_impl_parent_implementedSystem_port_0_cast <= Delay1No644_out;
Delay1No645_out_to_Subtract27_1_impl_parent_implementedSystem_port_1_cast <= Delay1No645_out;
   Subtract27_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract27_1_impl_out,
                 X => Delay1No644_out_to_Subtract27_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No645_out_to_Subtract27_1_impl_parent_implementedSystem_port_1_cast);

SharedReg760_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg760_out;
SharedReg406_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg406_out;
SharedReg7_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg7_out;
SharedReg761_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg761_out;
SharedReg384_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg384_out;
SharedReg527_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg527_out;
   MUX_Subtract27_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg760_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg406_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg7_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg761_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg384_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Subtract27_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_1_impl_0_out);

   Delay1No644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_1_impl_0_out,
                 Y => Delay1No644_out);

SharedReg790_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg790_out;
SharedReg440_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg440_out;
SharedReg23_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg791_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg791_out;
SharedReg627_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg226_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg226_out;
   MUX_Subtract27_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg790_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg440_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg23_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg791_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg226_out_to_MUX_Subtract27_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_1_impl_1_out);

   Delay1No645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_1_impl_1_out,
                 Y => Delay1No645_out);

Delay1No646_out_to_Subtract27_2_impl_parent_implementedSystem_port_0_cast <= Delay1No646_out;
Delay1No647_out_to_Subtract27_2_impl_parent_implementedSystem_port_1_cast <= Delay1No647_out;
   Subtract27_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract27_2_impl_out,
                 X => Delay1No646_out_to_Subtract27_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No647_out_to_Subtract27_2_impl_parent_implementedSystem_port_1_cast);

SharedReg615_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg615_out;
SharedReg685_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg685_out;
SharedReg251_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg251_out;
SharedReg6_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg6_out;
SharedReg763_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg763_out;
SharedReg358_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg358_out;
   MUX_Subtract27_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg615_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg685_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg251_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg763_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg358_out_to_MUX_Subtract27_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_2_impl_0_out);

   Delay1No646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_2_impl_0_out,
                 Y => Delay1No646_out);

SharedReg441_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg441_out;
SharedReg710_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg710_out;
SharedReg267_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg267_out;
SharedReg22_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
SharedReg793_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg793_out;
SharedReg648_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg648_out;
   MUX_Subtract27_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg441_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg710_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg267_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg793_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg648_out_to_MUX_Subtract27_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_2_impl_1_out);

   Delay1No647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_2_impl_1_out,
                 Y => Delay1No647_out);

Delay1No648_out_to_Subtract27_3_impl_parent_implementedSystem_port_0_cast <= Delay1No648_out;
Delay1No649_out_to_Subtract27_3_impl_parent_implementedSystem_port_1_cast <= Delay1No649_out;
   Subtract27_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract27_3_impl_out,
                 X => Delay1No648_out_to_Subtract27_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No649_out_to_Subtract27_3_impl_parent_implementedSystem_port_1_cast);

SharedReg238_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg238_out;
SharedReg535_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg535_out;
Delay3No218_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_3_cast <= Delay3No218_out;
SharedReg669_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg669_out;
SharedReg6_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg6_out;
SharedReg765_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg765_out;
   MUX_Subtract27_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg238_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg535_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No218_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg669_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg6_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg765_out_to_MUX_Subtract27_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_3_impl_0_out);

   Delay1No648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_3_impl_0_out,
                 Y => Delay1No648_out);

SharedReg536_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg536_out;
SharedReg236_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg236_out;
Delay3No223_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_3_cast <= Delay3No223_out;
SharedReg691_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg691_out;
SharedReg22_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg22_out;
SharedReg795_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg795_out;
   MUX_Subtract27_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg536_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg236_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No223_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg691_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg22_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg795_out_to_MUX_Subtract27_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_3_impl_1_out);

   Delay1No649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_3_impl_1_out,
                 Y => Delay1No649_out);

Delay1No650_out_to_Subtract27_4_impl_parent_implementedSystem_port_0_cast <= Delay1No650_out;
Delay1No651_out_to_Subtract27_4_impl_parent_implementedSystem_port_1_cast <= Delay1No651_out;
   Subtract27_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract27_4_impl_out,
                 X => Delay1No650_out_to_Subtract27_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No651_out_to_Subtract27_4_impl_parent_implementedSystem_port_1_cast);

SharedReg7_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg7_out;
SharedReg767_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg767_out;
SharedReg452_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg452_out;
SharedReg633_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg633_out;
SharedReg687_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg687_out;
SharedReg333_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg333_out;
   MUX_Subtract27_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg7_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg767_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg452_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg633_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg687_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg333_out_to_MUX_Subtract27_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_4_impl_0_out);

   Delay1No650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_4_impl_0_out,
                 Y => Delay1No650_out);

SharedReg23_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg23_out;
SharedReg797_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg797_out;
SharedReg756_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg756_out;
SharedReg393_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg393_out;
SharedReg714_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg714_out;
SharedReg396_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg396_out;
   MUX_Subtract27_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg23_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg797_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg756_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg393_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg714_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg396_out_to_MUX_Subtract27_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract27_4_impl_1_out);

   Delay1No651_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract27_4_impl_1_out,
                 Y => Delay1No651_out);

Delay1No652_out_to_Subtract42_0_impl_parent_implementedSystem_port_0_cast <= Delay1No652_out;
Delay1No653_out_to_Subtract42_0_impl_parent_implementedSystem_port_1_cast <= Delay1No653_out;
   Subtract42_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_0_impl_out,
                 X => Delay1No652_out_to_Subtract42_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No653_out_to_Subtract42_0_impl_parent_implementedSystem_port_1_cast);

SharedReg696_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg696_out;
SharedReg11_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg11_out;
SharedReg88_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg523_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg523_out;
SharedReg316_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg316_out;
SharedReg246_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg246_out;
   MUX_Subtract42_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg696_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg11_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg523_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg316_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg246_out_to_MUX_Subtract42_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_0_impl_0_out);

   Delay1No652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_0_impl_0_out,
                 Y => Delay1No652_out);

SharedReg586_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg586_out;
SharedReg27_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg27_out;
SharedReg523_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg523_out;
SharedReg277_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg277_out;
SharedReg636_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg636_out;
SharedReg119_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg119_out;
   MUX_Subtract42_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg586_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg523_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg277_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg636_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg119_out_to_MUX_Subtract42_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_0_impl_1_out);

   Delay1No653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_0_impl_1_out,
                 Y => Delay1No653_out);

Delay1No654_out_to_Subtract42_1_impl_parent_implementedSystem_port_0_cast <= Delay1No654_out;
Delay1No655_out_to_Subtract42_1_impl_parent_implementedSystem_port_1_cast <= Delay1No655_out;
   Subtract42_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_1_impl_out,
                 X => Delay1No654_out_to_Subtract42_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No655_out_to_Subtract42_1_impl_parent_implementedSystem_port_1_cast);

SharedReg228_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg228_out;
SharedReg698_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg698_out;
SharedReg11_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg92_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg92_out;
SharedReg406_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg406_out;
SharedReg174_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg174_out;
   MUX_Subtract42_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg228_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg698_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg11_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg406_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg174_out_to_MUX_Subtract42_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_1_impl_0_out);

   Delay1No654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_1_impl_0_out,
                 Y => Delay1No654_out);

SharedReg136_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg588_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg588_out;
SharedReg27_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg527_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg527_out;
SharedReg816_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg816_out;
SharedReg278_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg278_out;
   MUX_Subtract42_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg588_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg27_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg527_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg816_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg278_out_to_MUX_Subtract42_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_1_impl_1_out);

   Delay1No655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_1_impl_1_out,
                 Y => Delay1No655_out);

Delay1No656_out_to_Subtract42_2_impl_parent_implementedSystem_port_0_cast <= Delay1No656_out;
Delay1No657_out_to_Subtract42_2_impl_parent_implementedSystem_port_1_cast <= Delay1No657_out;
   Subtract42_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_2_impl_out,
                 X => Delay1No656_out_to_Subtract42_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No657_out_to_Subtract42_2_impl_parent_implementedSystem_port_1_cast);

SharedReg195_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg195_out;
SharedReg233_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg233_out;
SharedReg700_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg700_out;
SharedReg11_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg326_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg282_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg282_out;
   MUX_Subtract42_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg195_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg233_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg700_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg326_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg282_out_to_MUX_Subtract42_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_2_impl_0_out);

   Delay1No656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_2_impl_0_out,
                 Y => Delay1No656_out);

SharedReg281_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg281_out;
SharedReg139_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg590_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg590_out;
SharedReg27_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg27_out;
SharedReg409_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg409_out;
SharedReg533_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg533_out;
   MUX_Subtract42_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg281_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg590_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg27_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg409_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg533_out_to_MUX_Subtract42_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_2_impl_1_out);

   Delay1No657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_2_impl_1_out,
                 Y => Delay1No657_out);

Delay1No658_out_to_Subtract42_3_impl_parent_implementedSystem_port_0_cast <= Delay1No658_out;
Delay1No659_out_to_Subtract42_3_impl_parent_implementedSystem_port_1_cast <= Delay1No659_out;
   Subtract42_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_3_impl_out,
                 X => Delay1No658_out_to_Subtract42_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No659_out_to_Subtract42_3_impl_parent_implementedSystem_port_1_cast);

SharedReg535_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg535_out;
SharedReg205_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg254_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg254_out;
SharedReg702_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg702_out;
SharedReg12_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg544_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg544_out;
   MUX_Subtract42_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg535_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg254_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg702_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg544_out_to_MUX_Subtract42_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_3_impl_0_out);

   Delay1No658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_3_impl_0_out,
                 Y => Delay1No658_out);

SharedReg545_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg545_out;
SharedReg534_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg534_out;
SharedReg142_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg592_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg592_out;
SharedReg28_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg222_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg222_out;
   MUX_Subtract42_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg545_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg534_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg592_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg222_out_to_MUX_Subtract42_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_3_impl_1_out);

   Delay1No659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_3_impl_1_out,
                 Y => Delay1No659_out);

Delay1No660_out_to_Subtract42_4_impl_parent_implementedSystem_port_0_cast <= Delay1No660_out;
Delay1No661_out_to_Subtract42_4_impl_parent_implementedSystem_port_1_cast <= Delay1No661_out;
   Subtract42_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract42_4_impl_out,
                 X => Delay1No660_out_to_Subtract42_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No661_out_to_Subtract42_4_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg662_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg662_out;
SharedReg394_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg394_out;
SharedReg397_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg397_out;
SharedReg395_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg395_out;
SharedReg704_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg704_out;
   MUX_Subtract42_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg662_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg394_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg395_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg704_out_to_MUX_Subtract42_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_4_impl_0_out);

   Delay1No660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_4_impl_0_out,
                 Y => Delay1No660_out);

SharedReg27_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg477_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg477_out;
SharedReg737_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg737_out;
SharedReg451_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg451_out;
SharedReg473_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg473_out;
SharedReg594_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg594_out;
   MUX_Subtract42_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg477_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg737_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg451_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg473_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg594_out_to_MUX_Subtract42_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract42_4_impl_1_out);

   Delay1No661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract42_4_impl_1_out,
                 Y => Delay1No661_out);

Delay1No662_out_to_Add84_4_impl_parent_implementedSystem_port_0_cast <= Delay1No662_out;
Delay1No663_out_to_Add84_4_impl_parent_implementedSystem_port_1_cast <= Delay1No663_out;
   Add84_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add84_4_impl_out,
                 X => Delay1No662_out_to_Add84_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No663_out_to_Add84_4_impl_parent_implementedSystem_port_1_cast);

SharedReg787_out_to_MUX_Add84_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg787_out;
SharedReg776_out_to_MUX_Add84_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg776_out;
   MUX_Add84_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg787_out_to_MUX_Add84_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg776_out_to_MUX_Add84_4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add84_4_impl_0_LUT_out,
                 oMux => MUX_Add84_4_impl_0_out);

   Delay1No662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add84_4_impl_0_out,
                 Y => Delay1No662_out);

SharedReg796_out_to_MUX_Add84_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg796_out;
SharedReg786_out_to_MUX_Add84_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg786_out;
   MUX_Add84_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg796_out_to_MUX_Add84_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg786_out_to_MUX_Add84_4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add84_4_impl_1_LUT_out,
                 oMux => MUX_Add84_4_impl_1_out);

   Delay1No663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add84_4_impl_1_out,
                 Y => Delay1No663_out);

Delay1No664_out_to_Subtract44_0_impl_parent_implementedSystem_port_0_cast <= Delay1No664_out;
Delay1No665_out_to_Subtract44_0_impl_parent_implementedSystem_port_1_cast <= Delay1No665_out;
   Subtract44_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_0_impl_out,
                 X => Delay1No664_out_to_Subtract44_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No665_out_to_Subtract44_0_impl_parent_implementedSystem_port_1_cast);

SharedReg758_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg758_out;
SharedReg12_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg318_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg435_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg435_out;
SharedReg171_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg171_out;
SharedReg353_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg353_out;
   MUX_Subtract44_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg758_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg318_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg435_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg171_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg353_out_to_MUX_Subtract44_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_0_impl_0_out);

   Delay1No664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_0_impl_0_out,
                 Y => Delay1No664_out);

SharedReg674_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg674_out;
SharedReg28_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg435_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg435_out;
SharedReg813_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg813_out;
SharedReg274_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg274_out;
SharedReg600_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg600_out;
   MUX_Subtract44_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg674_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg435_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg813_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg274_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg600_out_to_MUX_Subtract44_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_0_impl_1_out);

   Delay1No665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_0_impl_1_out,
                 Y => Delay1No665_out);

Delay1No666_out_to_Subtract44_1_impl_parent_implementedSystem_port_0_cast <= Delay1No666_out;
Delay1No667_out_to_Subtract44_1_impl_parent_implementedSystem_port_1_cast <= Delay1No667_out;
   Subtract44_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_1_impl_out,
                 X => Delay1No666_out_to_Subtract44_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No667_out_to_Subtract44_1_impl_parent_implementedSystem_port_1_cast);

SharedReg386_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg386_out;
SharedReg760_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg760_out;
SharedReg12_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg322_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg322_out;
SharedReg527_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg527_out;
SharedReg355_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg355_out;
   MUX_Subtract44_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg386_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg760_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg12_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg322_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg527_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg355_out_to_MUX_Subtract44_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_1_impl_0_out);

   Delay1No666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_1_impl_0_out,
                 Y => Delay1No666_out);

SharedReg603_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg603_out;
SharedReg676_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg676_out;
SharedReg28_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg439_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg439_out;
SharedReg529_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg529_out;
SharedReg742_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg742_out;
   MUX_Subtract44_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg603_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg676_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg28_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg439_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg529_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg742_out_to_MUX_Subtract44_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_1_impl_1_out);

   Delay1No667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_1_impl_1_out,
                 Y => Delay1No667_out);

Delay1No668_out_to_Subtract44_2_impl_parent_implementedSystem_port_0_cast <= Delay1No668_out;
Delay1No669_out_to_Subtract44_2_impl_parent_implementedSystem_port_1_cast <= Delay1No669_out;
   Subtract44_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_2_impl_out,
                 X => Delay1No668_out_to_Subtract44_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No669_out_to_Subtract44_2_impl_parent_implementedSystem_port_1_cast);

SharedReg358_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg358_out;
SharedReg359_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg359_out;
SharedReg762_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg762_out;
SharedReg12_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg12_out;
SharedReg155_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg155_out;
SharedReg409_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg409_out;
   MUX_Subtract44_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg358_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg359_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg762_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg12_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg155_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg409_out_to_MUX_Subtract44_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_2_impl_0_out);

   Delay1No668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_2_impl_0_out,
                 Y => Delay1No668_out);

SharedReg803_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg803_out;
SharedReg615_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg615_out;
SharedReg678_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg678_out;
SharedReg28_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg28_out;
SharedReg218_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg218_out;
SharedReg839_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg839_out;
   MUX_Subtract44_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg803_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg615_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg678_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg28_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg218_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg839_out_to_MUX_Subtract44_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_2_impl_1_out);

   Delay1No669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_2_impl_1_out,
                 Y => Delay1No669_out);

Delay1No670_out_to_Subtract44_3_impl_parent_implementedSystem_port_0_cast <= Delay1No670_out;
Delay1No671_out_to_Subtract44_3_impl_parent_implementedSystem_port_1_cast <= Delay1No671_out;
   Subtract44_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_3_impl_out,
                 X => Delay1No670_out_to_Subtract44_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No671_out_to_Subtract44_3_impl_parent_implementedSystem_port_1_cast);

SharedReg412_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg412_out;
SharedReg361_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg361_out;
SharedReg521_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg521_out;
SharedReg764_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg764_out;
SharedReg13_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg447_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg447_out;
   MUX_Subtract44_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg412_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg361_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg521_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg764_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg447_out_to_MUX_Subtract44_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_3_impl_0_out);

   Delay1No670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_3_impl_0_out,
                 Y => Delay1No670_out);

SharedReg842_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg842_out;
SharedReg847_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg847_out;
SharedReg618_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg618_out;
SharedReg680_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg680_out;
SharedReg29_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg29_out;
SharedReg805_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg805_out;
   MUX_Subtract44_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg842_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg847_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg618_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg680_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg29_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg805_out_to_MUX_Subtract44_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_3_impl_1_out);

   Delay1No671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_3_impl_1_out,
                 Y => Delay1No671_out);

Delay1No672_out_to_Subtract44_4_impl_parent_implementedSystem_port_0_cast <= Delay1No672_out;
Delay1No673_out_to_Subtract44_4_impl_parent_implementedSystem_port_1_cast <= Delay1No673_out;
   Subtract44_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract44_4_impl_out,
                 X => Delay1No672_out_to_Subtract44_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No673_out_to_Subtract44_4_impl_parent_implementedSystem_port_1_cast);

SharedReg12_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg399_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg547_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg547_out;
SharedReg191_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg191_out;
SharedReg288_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg288_out;
SharedReg766_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg766_out;
   MUX_Subtract44_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg547_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg191_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg288_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg766_out_to_MUX_Subtract44_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_4_impl_0_out);

   Delay1No672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_4_impl_0_out,
                 Y => Delay1No672_out);

SharedReg28_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg28_out;
SharedReg394_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg394_out;
SharedReg290_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg477_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg477_out;
SharedReg103_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg103_out;
SharedReg682_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg682_out;
   MUX_Subtract44_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg28_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg394_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg290_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg477_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg103_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg682_out_to_MUX_Subtract44_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract44_4_impl_1_out);

   Delay1No673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract44_4_impl_1_out,
                 Y => Delay1No673_out);

Delay1No674_out_to_Subtract45_3_impl_parent_implementedSystem_port_0_cast <= Delay1No674_out;
Delay1No675_out_to_Subtract45_3_impl_parent_implementedSystem_port_1_cast <= Delay1No675_out;
   Subtract45_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract45_3_impl_out,
                 X => Delay1No674_out_to_Subtract45_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No675_out_to_Subtract45_3_impl_parent_implementedSystem_port_1_cast);

SharedReg361_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg361_out;
SharedReg618_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg618_out;
SharedReg686_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg686_out;
SharedReg269_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg269_out;
SharedReg7_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg7_out;
SharedReg362_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg362_out;
   MUX_Subtract45_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg361_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg618_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg686_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg269_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg7_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg362_out_to_MUX_Subtract45_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract45_3_impl_0_out);

   Delay1No674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_3_impl_0_out,
                 Y => Delay1No674_out);

SharedReg733_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg733_out;
SharedReg446_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg446_out;
SharedReg712_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg712_out;
SharedReg286_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg286_out;
SharedReg23_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg23_out;
SharedReg618_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg618_out;
   MUX_Subtract45_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg733_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg446_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg712_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg286_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg23_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg618_out_to_MUX_Subtract45_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract45_3_impl_1_out);

   Delay1No675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract45_3_impl_1_out,
                 Y => Delay1No675_out);

Delay1No676_out_to_Subtract46_0_impl_parent_implementedSystem_port_0_cast <= Delay1No676_out;
Delay1No677_out_to_Subtract46_0_impl_parent_implementedSystem_port_1_cast <= Delay1No677_out;
   Subtract46_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_0_impl_out,
                 X => Delay1No676_out_to_Subtract46_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No677_out_to_Subtract46_0_impl_parent_implementedSystem_port_1_cast);

SharedReg778_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg778_out;
SharedReg13_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg540_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg540_out;
SharedReg539_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg539_out;
SharedReg351_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg621_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg621_out;
   MUX_Subtract46_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg778_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg540_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg539_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg621_out_to_MUX_Subtract46_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_0_impl_0_out);

   Delay1No676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_0_impl_0_out,
                 Y => Delay1No676_out);

Delay3No235_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_1_cast <= Delay3No235_out;
SharedReg29_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg224_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg224_out;
SharedReg525_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg525_out;
SharedReg738_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg738_out;
SharedReg319_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg319_out;
   MUX_Subtract46_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No235_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg224_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg525_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg738_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg319_out_to_MUX_Subtract46_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_0_impl_1_out);

   Delay1No677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_0_impl_1_out,
                 Y => Delay1No677_out);

Delay1No678_out_to_Subtract46_1_impl_parent_implementedSystem_port_0_cast <= Delay1No678_out;
Delay1No679_out_to_Subtract46_1_impl_parent_implementedSystem_port_1_cast <= Delay1No679_out;
   Subtract46_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_1_impl_out,
                 X => Delay1No678_out_to_Subtract46_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No679_out_to_Subtract46_1_impl_parent_implementedSystem_port_1_cast);

SharedReg625_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg625_out;
SharedReg780_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg780_out;
SharedReg13_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg150_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg150_out;
SharedReg439_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg439_out;
SharedReg214_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg214_out;
   MUX_Subtract46_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg625_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg780_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg13_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg150_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg439_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg214_out_to_MUX_Subtract46_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_1_impl_0_out);

   Delay1No678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_1_impl_0_out,
                 Y => Delay1No678_out);

SharedReg323_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg323_out;
Delay3No236_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_2_cast <= Delay3No236_out;
SharedReg29_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg227_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg227_out;
SharedReg835_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg526_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg526_out;
   MUX_Subtract46_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg323_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No236_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg29_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg227_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg526_out_to_MUX_Subtract46_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_1_impl_1_out);

   Delay1No679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_1_impl_1_out,
                 Y => Delay1No679_out);

Delay1No680_out_to_Subtract46_2_impl_parent_implementedSystem_port_0_cast <= Delay1No680_out;
Delay1No681_out_to_Subtract46_2_impl_parent_implementedSystem_port_1_cast <= Delay1No681_out;
   Subtract46_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_2_impl_out,
                 X => Delay1No680_out_to_Subtract46_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No681_out_to_Subtract46_2_impl_parent_implementedSystem_port_1_cast);

SharedReg218_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg218_out;
SharedReg646_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg646_out;
SharedReg782_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg782_out;
SharedReg13_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg13_out;
SharedReg615_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg615_out;
SharedReg531_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg531_out;
   MUX_Subtract46_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg218_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg646_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg782_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg13_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg615_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg531_out_to_MUX_Subtract46_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_2_impl_0_out);

   Delay1No680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_2_impl_0_out,
                 Y => Delay1No680_out);

SharedReg530_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg530_out;
SharedReg327_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg327_out;
Delay3No237_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_3_cast <= Delay3No237_out;
SharedReg29_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg29_out;
SharedReg804_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg804_out;
SharedReg157_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg157_out;
   MUX_Subtract46_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg530_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg327_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No237_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg29_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg804_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg157_out_to_MUX_Subtract46_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_2_impl_1_out);

   Delay1No681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_2_impl_1_out,
                 Y => Delay1No681_out);

Delay1No682_out_to_Subtract46_3_impl_parent_implementedSystem_port_0_cast <= Delay1No682_out;
Delay1No683_out_to_Subtract46_3_impl_parent_implementedSystem_port_1_cast <= Delay1No683_out;
   Subtract46_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_3_impl_out,
                 X => Delay1No682_out_to_Subtract46_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No683_out_to_Subtract46_3_impl_parent_implementedSystem_port_1_cast);

SharedReg543_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg543_out;
SharedReg237_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg237_out;
SharedReg731_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg731_out;
SharedReg784_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg784_out;
SharedReg14_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg14_out;
SharedReg253_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg253_out;
   MUX_Subtract46_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg543_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg237_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg731_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg784_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg14_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg253_out_to_MUX_Subtract46_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_3_impl_0_out);

   Delay1No682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_3_impl_0_out,
                 Y => Delay1No682_out);

SharedReg48_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg542_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg542_out;
SharedReg331_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg331_out;
Delay3No238_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_4_cast <= Delay3No238_out;
SharedReg30_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg543_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg543_out;
   MUX_Subtract46_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg542_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg331_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No238_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg543_out_to_MUX_Subtract46_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_3_impl_1_out);

   Delay1No683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_3_impl_1_out,
                 Y => Delay1No683_out);

Delay1No684_out_to_Subtract46_4_impl_parent_implementedSystem_port_0_cast <= Delay1No684_out;
Delay1No685_out_to_Subtract46_4_impl_parent_implementedSystem_port_1_cast <= Delay1No685_out;
   Subtract46_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_4_impl_out,
                 X => Delay1No684_out_to_Subtract46_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No685_out_to_Subtract46_4_impl_parent_implementedSystem_port_1_cast);

SharedReg13_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg13_out;
SharedReg548_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg548_out;
SharedReg451_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg451_out;
SharedReg332_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg332_out;
SharedReg475_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg475_out;
SharedReg786_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg786_out;
   MUX_Subtract46_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg13_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg548_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg451_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg332_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg475_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg786_out_to_MUX_Subtract46_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_4_impl_0_out);

   Delay1No684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_4_impl_0_out,
                 Y => Delay1No684_out);

SharedReg29_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg29_out;
SharedReg242_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg242_out;
SharedReg826_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg826_out;
SharedReg734_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg734_out;
SharedReg596_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg596_out;
Delay3No239_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_6_cast <= Delay3No239_out;
   MUX_Subtract46_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg242_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg826_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg734_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg596_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay3No239_out_to_MUX_Subtract46_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract46_4_impl_1_out);

   Delay1No685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_4_impl_1_out,
                 Y => Delay1No685_out);

Delay1No686_out_to_Subtract47_2_impl_parent_implementedSystem_port_0_cast <= Delay1No686_out;
Delay1No687_out_to_Subtract47_2_impl_parent_implementedSystem_port_1_cast <= Delay1No687_out;
   Subtract47_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract47_2_impl_out,
                 X => Delay1No686_out_to_Subtract47_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No687_out_to_Subtract47_2_impl_parent_implementedSystem_port_1_cast);

SharedReg531_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg531_out;
SharedReg762_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg762_out;
SharedReg409_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg409_out;
SharedReg7_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg7_out;
SharedReg389_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg389_out;
SharedReg251_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg251_out;
   MUX_Subtract47_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg531_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg762_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg409_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg7_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg389_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg251_out_to_MUX_Subtract47_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract47_2_impl_0_out);

   Delay1No686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_2_impl_0_out,
                 Y => Delay1No686_out);

SharedReg231_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg231_out;
SharedReg792_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg445_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg445_out;
SharedReg23_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
SharedReg629_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg629_out;
SharedReg235_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg235_out;
   MUX_Subtract47_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg231_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg445_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg23_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg629_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg235_out_to_MUX_Subtract47_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract47_2_impl_1_out);

   Delay1No687_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_2_impl_1_out,
                 Y => Delay1No687_out);

Delay1No688_out_to_Subtract47_3_impl_parent_implementedSystem_port_0_cast <= Delay1No688_out;
Delay1No689_out_to_Subtract47_3_impl_parent_implementedSystem_port_1_cast <= Delay1No689_out;
   Subtract47_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract47_3_impl_out,
                 X => Delay1No688_out_to_Subtract47_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No689_out_to_Subtract47_3_impl_parent_implementedSystem_port_1_cast);

SharedReg269_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg269_out;
SharedReg543_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg543_out;
SharedReg764_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg764_out;
SharedReg412_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg412_out;
SharedReg8_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg8_out;
SharedReg536_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg536_out;
   MUX_Subtract47_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg269_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg543_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg764_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg412_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg8_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg536_out_to_MUX_Subtract47_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract47_3_impl_0_out);

   Delay1No688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_3_impl_0_out,
                 Y => Delay1No688_out);

SharedReg256_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg252_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg252_out;
SharedReg794_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg794_out;
SharedReg449_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg449_out;
SharedReg24_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg24_out;
SharedReg269_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg269_out;
   MUX_Subtract47_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg794_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg449_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg24_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg269_out_to_MUX_Subtract47_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract47_3_impl_1_out);

   Delay1No689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_3_impl_1_out,
                 Y => Delay1No689_out);

Delay1No690_out_to_Subtract47_4_impl_parent_implementedSystem_port_0_cast <= Delay1No690_out;
Delay1No691_out_to_Subtract47_4_impl_parent_implementedSystem_port_1_cast <= Delay1No691_out;
   Subtract47_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract47_4_impl_out,
                 X => Delay1No690_out_to_Subtract47_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No691_out_to_Subtract47_4_impl_parent_implementedSystem_port_1_cast);

SharedReg8_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg474_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg474_out;
Delay3No134_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_3_cast <= Delay3No134_out;
SharedReg661_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg661_out;
SharedReg766_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg766_out;
SharedReg131_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg131_out;
   MUX_Subtract47_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg474_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No134_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg661_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg766_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg131_out_to_MUX_Subtract47_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract47_4_impl_0_out);

   Delay1No690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_4_impl_0_out,
                 Y => Delay1No690_out);

SharedReg24_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg633_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg633_out;
SharedReg548_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg548_out;
SharedReg241_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg241_out;
SharedReg796_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg796_out;
SharedReg147_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
   MUX_Subtract47_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg633_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg548_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg796_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg147_out_to_MUX_Subtract47_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract47_4_impl_1_out);

   Delay1No691_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_4_impl_1_out,
                 Y => Delay1No691_out);

Delay1No692_out_to_Subtract52_0_impl_parent_implementedSystem_port_0_cast <= Delay1No692_out;
Delay1No693_out_to_Subtract52_0_impl_parent_implementedSystem_port_1_cast <= Delay1No693_out;
   Subtract52_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract52_0_impl_out,
                 X => Delay1No692_out_to_Subtract52_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No693_out_to_Subtract52_0_impl_parent_implementedSystem_port_1_cast);

SharedReg162_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg162_out;
SharedReg8_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg352_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg352_out;
SharedReg317_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg317_out;
SharedReg539_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg539_out;
SharedReg436_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg436_out;
   MUX_Subtract52_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg162_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg352_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg317_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg539_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg436_out_to_MUX_Subtract52_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_0_impl_0_out);

   Delay1No692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_0_impl_0_out,
                 Y => Delay1No692_out);

SharedReg173_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg173_out;
SharedReg24_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg621_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg621_out;
SharedReg623_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg623_out;
SharedReg223_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg223_out;
SharedReg849_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg849_out;
   MUX_Subtract52_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg173_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg621_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg623_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg223_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg849_out_to_MUX_Subtract52_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_0_impl_1_out);

   Delay1No693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_0_impl_1_out,
                 Y => Delay1No693_out);

Delay1No694_out_to_Subtract52_1_impl_parent_implementedSystem_port_0_cast <= Delay1No694_out;
Delay1No695_out_to_Subtract52_1_impl_parent_implementedSystem_port_1_cast <= Delay1No695_out;
   Subtract52_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract52_1_impl_out,
                 X => Delay1No694_out_to_Subtract52_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No695_out_to_Subtract52_1_impl_parent_implementedSystem_port_1_cast);

SharedReg407_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg407_out;
SharedReg165_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg8_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg385_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg385_out;
SharedReg262_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg262_out;
SharedReg383_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg383_out;
   MUX_Subtract52_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg407_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg8_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg385_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg262_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg383_out_to_MUX_Subtract52_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_1_impl_0_out);

   Delay1No694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_1_impl_0_out,
                 Y => Delay1No694_out);

SharedReg851_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg851_out;
SharedReg176_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg176_out;
SharedReg24_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg625_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg625_out;
SharedReg230_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg230_out;
SharedReg321_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg321_out;
   MUX_Subtract52_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg851_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg176_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg625_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg230_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg321_out_to_MUX_Subtract52_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_1_impl_1_out);

   Delay1No695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_1_impl_1_out,
                 Y => Delay1No695_out);

Delay1No696_out_to_Subtract52_2_impl_parent_implementedSystem_port_0_cast <= Delay1No696_out;
Delay1No697_out_to_Subtract52_2_impl_parent_implementedSystem_port_1_cast <= Delay1No697_out;
   Subtract52_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract52_2_impl_out,
                 X => Delay1No696_out_to_Subtract52_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No697_out_to_Subtract52_2_impl_parent_implementedSystem_port_1_cast);

SharedReg387_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg387_out;
SharedReg410_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg410_out;
SharedReg178_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg178_out;
SharedReg8_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg8_out;
SharedReg532_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg532_out;
SharedReg388_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg388_out;
   MUX_Subtract52_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg387_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg410_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg178_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg8_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg532_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg388_out_to_MUX_Subtract52_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_2_impl_0_out);

   Delay1No696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_2_impl_0_out,
                 Y => Delay1No696_out);

SharedReg325_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg325_out;
SharedReg853_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg853_out;
SharedReg198_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg24_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg24_out;
SharedReg265_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg748_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg748_out;
   MUX_Subtract52_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg325_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg853_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg198_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg24_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg748_out_to_MUX_Subtract52_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_2_impl_1_out);

   Delay1No697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_2_impl_1_out,
                 Y => Delay1No697_out);

Delay1No698_out_to_Subtract52_3_impl_parent_implementedSystem_port_0_cast <= Delay1No698_out;
Delay1No699_out_to_Subtract52_3_impl_parent_implementedSystem_port_1_cast <= Delay1No699_out;
   Subtract52_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract52_3_impl_out,
                 X => Delay1No698_out_to_Subtract52_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No699_out_to_Subtract52_3_impl_parent_implementedSystem_port_1_cast);

SharedReg391_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg390_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg390_out;
SharedReg413_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg183_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg183_out;
SharedReg9_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg9_out;
SharedReg330_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg330_out;
   MUX_Subtract52_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg390_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg413_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg183_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg9_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg330_out_to_MUX_Subtract52_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_3_impl_0_out);

   Delay1No698_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_3_impl_0_out,
                 Y => Delay1No698_out);

SharedReg807_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg807_out;
SharedReg329_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg329_out;
SharedReg855_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg855_out;
SharedReg208_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg208_out;
SharedReg25_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg25_out;
SharedReg731_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg731_out;
   MUX_Subtract52_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg807_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg329_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg855_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg208_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg25_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg731_out_to_MUX_Subtract52_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_3_impl_1_out);

   Delay1No699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_3_impl_1_out,
                 Y => Delay1No699_out);

Delay1No700_out_to_Subtract52_4_impl_parent_implementedSystem_port_0_cast <= Delay1No700_out;
Delay1No701_out_to_Subtract52_4_impl_parent_implementedSystem_port_1_cast <= Delay1No701_out;
   Subtract52_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract52_4_impl_out,
                 X => Delay1No700_out_to_Subtract52_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No701_out_to_Subtract52_4_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg478_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg478_out;
SharedReg333_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg333_out;
SharedReg656_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg656_out;
SharedReg597_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg597_out;
SharedReg451_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg451_out;
   MUX_Subtract52_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg478_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg333_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg656_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg597_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg451_out_to_MUX_Subtract52_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_4_impl_0_out);

   Delay1No700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_4_impl_0_out,
                 Y => Delay1No700_out);

SharedReg25_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg287_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg287_out;
SharedReg635_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg635_out;
SharedReg450_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg450_out;
SharedReg856_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg856_out;
SharedReg598_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg598_out;
   MUX_Subtract52_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg287_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg635_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg450_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg856_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg598_out_to_MUX_Subtract52_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract52_4_impl_1_out);

   Delay1No701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract52_4_impl_1_out,
                 Y => Delay1No701_out);

Delay1No702_out_to_Subtract112_0_impl_parent_implementedSystem_port_0_cast <= Delay1No702_out;
Delay1No703_out_to_Subtract112_0_impl_parent_implementedSystem_port_1_cast <= Delay1No703_out;
   Subtract112_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract112_0_impl_out,
                 X => Delay1No702_out_to_Subtract112_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No703_out_to_Subtract112_0_impl_parent_implementedSystem_port_1_cast);

SharedReg600_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg600_out;
SharedReg9_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg524_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg524_out;
SharedReg275_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg275_out;
SharedReg350_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg350_out;
SharedReg276_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg276_out;
   MUX_Subtract112_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg600_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg524_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg275_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg350_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg276_out_to_MUX_Subtract112_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_0_impl_0_out);

   Delay1No702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_0_impl_0_out,
                 Y => Delay1No702_out);

SharedReg609_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg609_out;
SharedReg25_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
SharedReg275_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg275_out;
SharedReg225_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg225_out;
SharedReg403_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg403_out;
SharedReg86_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg86_out;
   MUX_Subtract112_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg609_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg275_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg225_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg403_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg86_out_to_MUX_Subtract112_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_0_impl_1_out);

   Delay1No703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_0_impl_1_out,
                 Y => Delay1No703_out);

Delay1No704_out_to_Subtract112_1_impl_parent_implementedSystem_port_0_cast <= Delay1No704_out;
Delay1No705_out_to_Subtract112_1_impl_parent_implementedSystem_port_1_cast <= Delay1No705_out;
   Subtract112_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract112_1_impl_out,
                 X => Delay1No704_out_to_Subtract112_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No705_out_to_Subtract112_1_impl_parent_implementedSystem_port_1_cast);

SharedReg263_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg263_out;
SharedReg603_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg603_out;
SharedReg9_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg528_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg528_out;
SharedReg321_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg321_out;
SharedReg199_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg199_out;
   MUX_Subtract112_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg263_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg603_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg528_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg321_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg199_out_to_MUX_Subtract112_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_1_impl_0_out);

   Delay1No704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_1_impl_0_out,
                 Y => Delay1No704_out);

SharedReg90_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg613_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg613_out;
SharedReg25_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg279_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg279_out;
SharedReg725_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg725_out;
SharedReg248_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg248_out;
   MUX_Subtract112_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg613_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg25_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg279_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg725_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg248_out_to_MUX_Subtract112_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_1_impl_1_out);

   Delay1No705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_1_impl_1_out,
                 Y => Delay1No705_out);

Delay1No706_out_to_Subtract112_2_impl_parent_implementedSystem_port_0_cast <= Delay1No706_out;
Delay1No707_out_to_Subtract112_2_impl_parent_implementedSystem_port_1_cast <= Delay1No707_out;
   Subtract112_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract112_2_impl_out,
                 X => Delay1No706_out_to_Subtract112_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No707_out_to_Subtract112_2_impl_parent_implementedSystem_port_1_cast);

SharedReg202_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg202_out;
SharedReg266_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg266_out;
SharedReg615_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg615_out;
SharedReg9_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg9_out;
SharedReg410_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg410_out;
SharedReg265_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg265_out;
   MUX_Subtract112_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg202_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg266_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg615_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg9_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg410_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg265_out_to_MUX_Subtract112_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_2_impl_0_out);

   Delay1No706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_2_impl_0_out,
                 Y => Delay1No706_out);

SharedReg251_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg251_out;
SharedReg41_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg631_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg631_out;
SharedReg25_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
SharedReg727_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg727_out;
SharedReg283_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg283_out;
   MUX_Subtract112_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg251_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg631_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg727_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg283_out_to_MUX_Subtract112_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_2_impl_1_out);

   Delay1No707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_2_impl_1_out,
                 Y => Delay1No707_out);

Delay1No708_out_to_Subtract112_3_impl_parent_implementedSystem_port_0_cast <= Delay1No708_out;
Delay1No709_out_to_Subtract112_3_impl_parent_implementedSystem_port_1_cast <= Delay1No709_out;
   Subtract112_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract112_3_impl_out,
                 X => Delay1No708_out_to_Subtract112_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No709_out_to_Subtract112_3_impl_parent_implementedSystem_port_1_cast);

SharedReg284_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg284_out;
SharedReg221_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg221_out;
SharedReg285_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg285_out;
SharedReg618_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg618_out;
SharedReg10_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg10_out;
SharedReg47_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg47_out;
   MUX_Subtract112_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg284_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg285_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg618_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg10_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg47_out_to_MUX_Subtract112_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_3_impl_0_out);

   Delay1No708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_3_impl_0_out,
                 Y => Delay1No708_out);

SharedReg537_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg537_out;
SharedReg269_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg269_out;
SharedReg60_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg60_out;
SharedReg654_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg654_out;
SharedReg26_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg26_out;
SharedReg284_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg284_out;
   MUX_Subtract112_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg537_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg269_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg60_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg654_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg26_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg284_out_to_MUX_Subtract112_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_3_impl_1_out);

   Delay1No709_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_3_impl_1_out,
                 Y => Delay1No709_out);

Delay1No710_out_to_Subtract112_4_impl_parent_implementedSystem_port_0_cast <= Delay1No710_out;
Delay1No711_out_to_Subtract112_4_impl_parent_implementedSystem_port_1_cast <= Delay1No711_out;
   Subtract112_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract112_4_impl_out,
                 X => Delay1No710_out_to_Subtract112_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No711_out_to_Subtract112_4_impl_parent_implementedSystem_port_1_cast);

SharedReg10_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg334_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg334_out;
SharedReg477_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg477_out;
SharedReg827_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg827_out;
SharedReg548_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg186_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg186_out;
   MUX_Subtract112_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg334_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg477_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg827_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg186_out_to_MUX_Subtract112_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_4_impl_0_out);

   Delay1No710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_4_impl_0_out,
                 Y => Delay1No710_out);

SharedReg26_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg735_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg735_out;
SharedReg243_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg243_out;
SharedReg257_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg257_out;
SharedReg660_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg660_out;
SharedReg194_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg194_out;
   MUX_Subtract112_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg735_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg243_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg257_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg660_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg194_out_to_MUX_Subtract112_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract112_4_impl_1_out);

   Delay1No711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract112_4_impl_1_out,
                 Y => Delay1No711_out);

Delay1No712_out_to_Subtract56_0_impl_parent_implementedSystem_port_0_cast <= Delay1No712_out;
Delay1No713_out_to_Subtract56_0_impl_parent_implementedSystem_port_1_cast <= Delay1No713_out;
   Subtract56_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract56_0_impl_out,
                 X => Delay1No712_out_to_Subtract56_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No713_out_to_Subtract56_0_impl_parent_implementedSystem_port_1_cast);

SharedReg189_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg10_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg404_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg404_out;
SharedReg403_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg403_out;
SharedReg188_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg188_out;
SharedReg318_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg318_out;
   MUX_Subtract56_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg404_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg403_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg188_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg318_out_to_MUX_Subtract56_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_0_impl_0_out);

   Delay1No712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_0_impl_0_out,
                 Y => Delay1No712_out);

SharedReg212_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg212_out;
SharedReg26_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg717_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg717_out;
SharedReg720_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg720_out;
SharedReg259_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg259_out;
SharedReg350_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg350_out;
   MUX_Subtract56_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg212_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg717_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg720_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg259_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg350_out_to_MUX_Subtract56_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_0_impl_1_out);

   Delay1No713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_0_impl_1_out,
                 Y => Delay1No713_out);

Delay1No714_out_to_Subtract56_1_impl_parent_implementedSystem_port_0_cast <= Delay1No714_out;
Delay1No715_out_to_Subtract56_1_impl_parent_implementedSystem_port_1_cast <= Delay1No715_out;
   Subtract56_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract56_1_impl_out,
                 X => Delay1No714_out_to_Subtract56_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No715_out_to_Subtract56_1_impl_parent_implementedSystem_port_1_cast);

SharedReg385_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg385_out;
SharedReg200_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg200_out;
SharedReg10_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg10_out;
SharedReg407_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg279_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg279_out;
SharedReg320_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg320_out;
   MUX_Subtract56_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg385_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg200_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg10_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg279_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg320_out_to_MUX_Subtract56_1_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_1_impl_0_out);

   Delay1No714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_1_impl_0_out,
                 Y => Delay1No714_out);

SharedReg383_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg383_out;
SharedReg216_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg216_out;
SharedReg26_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg722_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg280_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg280_out;
SharedReg640_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg640_out;
   MUX_Subtract56_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg383_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg216_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg26_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg280_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg640_out_to_MUX_Subtract56_1_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_1_impl_1_out);

   Delay1No715_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_1_impl_1_out,
                 Y => Delay1No715_out);

Delay1No716_out_to_Subtract56_2_impl_parent_implementedSystem_port_0_cast <= Delay1No716_out;
Delay1No717_out_to_Subtract56_2_impl_parent_implementedSystem_port_1_cast <= Delay1No717_out;
   Subtract56_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract56_2_impl_out,
                 X => Delay1No716_out_to_Subtract56_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No717_out_to_Subtract56_2_impl_parent_implementedSystem_port_1_cast);

SharedReg324_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg324_out;
SharedReg389_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg203_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg203_out;
SharedReg10_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg10_out;
SharedReg43_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg43_out;
SharedReg325_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg325_out;
   MUX_Subtract56_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg324_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg203_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg10_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg43_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg325_out_to_MUX_Subtract56_2_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_2_impl_0_out);

   Delay1No716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_2_impl_0_out,
                 Y => Delay1No716_out);

SharedReg726_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg726_out;
SharedReg387_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg387_out;
SharedReg220_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg26_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg282_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg282_out;
SharedReg819_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg819_out;
   MUX_Subtract56_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg726_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg387_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg220_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg282_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg819_out_to_MUX_Subtract56_2_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_2_impl_1_out);

   Delay1No717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_2_impl_1_out,
                 Y => Delay1No717_out);

Delay1No718_out_to_Subtract56_3_impl_parent_implementedSystem_port_0_cast <= Delay1No718_out;
Delay1No719_out_to_Subtract56_3_impl_parent_implementedSystem_port_1_cast <= Delay1No719_out;
   Subtract56_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract56_3_impl_out,
                 X => Delay1No718_out_to_Subtract56_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No719_out_to_Subtract56_3_impl_parent_implementedSystem_port_1_cast);

SharedReg329_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg329_out;
SharedReg328_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg328_out;
SharedReg392_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg222_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg222_out;
SharedReg11_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg11_out;
SharedReg392_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg392_out;
   MUX_Subtract56_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg329_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg328_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg222_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg11_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg392_out_to_MUX_Subtract56_3_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_3_impl_0_out);

   Delay1No718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_3_impl_0_out,
                 Y => Delay1No718_out);

SharedReg823_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg823_out;
SharedReg749_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg749_out;
SharedReg390_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg240_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg240_out;
SharedReg27_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg27_out;
SharedReg329_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg329_out;
   MUX_Subtract56_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg823_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg749_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg240_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg27_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg329_out_to_MUX_Subtract56_3_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract56_3_impl_1_out);

   Delay1No719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract56_3_impl_1_out,
                 Y => Delay1No719_out);

Delay1No720_out_to_Subtract60_0_impl_parent_implementedSystem_port_0_cast <= Delay1No720_out;
Delay1No721_out_to_Subtract60_0_impl_parent_implementedSystem_port_1_cast <= Delay1No721_out;
   Subtract60_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract60_0_impl_out,
                 X => Delay1No720_out_to_Subtract60_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No721_out_to_Subtract60_0_impl_parent_implementedSystem_port_1_cast);

SharedReg638_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg638_out;
SharedReg14_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg607_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg607_out;
SharedReg600_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg600_out;
SharedReg224_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg224_out;
SharedReg259_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg259_out;
   MUX_Subtract60_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg638_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg607_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg600_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg224_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg259_out_to_MUX_Subtract60_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract60_0_impl_0_out);

   Delay1No720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract60_0_impl_0_out,
                 Y => Delay1No720_out);

SharedReg353_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg30_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg799_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg799_out;
SharedReg831_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg831_out;
SharedReg522_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg522_out;
SharedReg135_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg135_out;
   MUX_Subtract60_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg799_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg831_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg522_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg135_out_to_MUX_Subtract60_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract60_0_impl_1_out);

   Delay1No721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract60_0_impl_1_out,
                 Y => Delay1No721_out);

Delay1No722_out_to_Subtract60_4_impl_parent_implementedSystem_port_0_cast <= Delay1No722_out;
Delay1No723_out_to_Subtract60_4_impl_parent_implementedSystem_port_1_cast <= Delay1No723_out;
   Subtract60_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract60_4_impl_out,
                 X => Delay1No722_out_to_Subtract60_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No723_out_to_Subtract60_4_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg596_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg596_out;
SharedReg661_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg661_out;
SharedReg185_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg185_out;
SharedReg656_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg656_out;
SharedReg658_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg658_out;
   MUX_Subtract60_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg596_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg661_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg185_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg656_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg658_out_to_MUX_Subtract60_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract60_4_impl_0_out);

   Delay1No722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract60_4_impl_0_out,
                 Y => Delay1No722_out);

SharedReg30_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg30_out;
SharedReg809_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg809_out;
SharedReg479_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg479_out;
SharedReg476_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg476_out;
SharedReg401_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg401_out;
SharedReg400_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg400_out;
   MUX_Subtract60_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg30_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg809_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg479_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg476_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg401_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Subtract60_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract60_4_impl_1_out);

   Delay1No723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract60_4_impl_1_out,
                 Y => Delay1No723_out);

Delay1No724_out_to_Subtract126_4_impl_parent_implementedSystem_port_0_cast <= Delay1No724_out;
Delay1No725_out_to_Subtract126_4_impl_parent_implementedSystem_port_1_cast <= Delay1No725_out;
   Subtract126_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract126_4_impl_out,
                 X => Delay1No724_out_to_Subtract126_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No725_out_to_Subtract126_4_impl_parent_implementedSystem_port_1_cast);

SharedReg15_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg15_out;
SharedReg271_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg271_out;
SharedReg596_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg596_out;
SharedReg333_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg333_out;
SharedReg287_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg287_out;
SharedReg756_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg756_out;
   MUX_Subtract126_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg271_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg596_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg333_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg287_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg756_out_to_MUX_Subtract126_4_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract126_4_impl_0_out);

   Delay1No724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract126_4_impl_0_out,
                 Y => Delay1No724_out);

SharedReg31_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg31_out;
SharedReg661_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg661_out;
SharedReg846_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg846_out;
SharedReg808_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg118_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg118_out;
Delay8No54_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_6_cast <= Delay8No54_out;
   MUX_Subtract126_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg31_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg661_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg846_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg118_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay8No54_out_to_MUX_Subtract126_4_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => ModCount61_out,
                 oMux => MUX_Subtract126_4_impl_1_out);

   Delay1No725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract126_4_impl_1_out,
                 Y => Delay1No725_out);

Delay1No726_out_to_Subtract135_4_impl_parent_implementedSystem_port_0_cast <= Delay1No726_out;
Delay1No727_out_to_Subtract135_4_impl_parent_implementedSystem_port_1_cast <= Delay1No727_out;
   Subtract135_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract135_4_impl_out,
                 X => Delay1No726_out_to_Subtract135_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No727_out_to_Subtract135_4_impl_parent_implementedSystem_port_1_cast);

SharedReg271_out_to_MUX_Subtract135_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg827_out_to_MUX_Subtract135_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg827_out;
   MUX_Subtract135_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Subtract135_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg827_out_to_MUX_Subtract135_4_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract135_4_impl_0_LUT_out,
                 oMux => MUX_Subtract135_4_impl_0_out);

   Delay1No726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract135_4_impl_0_out,
                 Y => Delay1No726_out);

SharedReg549_out_to_MUX_Subtract135_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg549_out;
SharedReg546_out_to_MUX_Subtract135_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg546_out;
   MUX_Subtract135_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg549_out_to_MUX_Subtract135_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg546_out_to_MUX_Subtract135_4_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract135_4_impl_1_LUT_out,
                 oMux => MUX_Subtract135_4_impl_1_out);

   Delay1No727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract135_4_impl_1_out,
                 Y => Delay1No727_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay3No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => Delay3No30_out);

   Delay3No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => Delay3No31_out);

   Delay3No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => Delay3No32_out);

   Delay3No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => Delay3No33_out);

   Delay3No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => Delay3No34_out);

   Delay3No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => Delay3No35_out);

   Delay3No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => Delay3No36_out);

   Delay3No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => Delay3No37_out);

   Delay3No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => Delay3No38_out);

   Delay3No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => Delay3No39_out);

   Delay2No320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => Delay2No320_out);

   Delay2No321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => Delay2No321_out);

   Delay2No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => Delay2No322_out);

   Delay2No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => Delay2No323_out);

   Delay2No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => Delay2No324_out);

   Delay2No325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => Delay2No325_out);

   Delay2No326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => Delay2No326_out);

   Delay2No327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => Delay2No327_out);

   Delay2No328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => Delay2No328_out);

   Delay2No329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => Delay2No329_out);

   Delay3No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => Delay3No134_out);

   Delay3No145_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => Delay3No145_out);

   Delay3No146_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => Delay3No146_out);

   Delay3No147_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => Delay3No147_out);

   Delay3No148_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => Delay3No148_out);

   Delay3No149_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => Delay3No149_out);

   Delay3No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => Delay3No150_out);

   Delay3No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => Delay3No151_out);

   Delay3No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => Delay3No152_out);

   Delay3No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => Delay3No153_out);

   Delay3No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => Delay3No154_out);

   Delay4No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => Delay4No40_out);

   Delay4No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay4No46_out);

   Delay3No195_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => Delay3No195_out);

   Delay3No196_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => Delay3No196_out);

   Delay3No197_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => Delay3No197_out);

   Delay3No198_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => Delay3No198_out);

   Delay3No199_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => Delay3No199_out);

   Delay3No200_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => Delay3No200_out);

   Delay3No201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => Delay3No201_out);

   Delay3No202_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => Delay3No202_out);

   Delay3No203_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => Delay3No203_out);

   Delay3No204_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => Delay3No204_out);

   Delay3No205_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => Delay3No205_out);

   Delay3No206_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => Delay3No206_out);

   Delay3No207_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => Delay3No207_out);

   Delay3No208_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => Delay3No208_out);

   Delay3No209_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => Delay3No209_out);

   Delay3No210_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => Delay3No210_out);

   Delay3No211_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => Delay3No211_out);

   Delay3No212_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => Delay3No212_out);

   Delay3No213_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => Delay3No213_out);

   Delay3No214_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => Delay3No214_out);

   Delay4No50_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => Delay4No50_out);

   Delay4No51_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => Delay4No51_out);

   Delay4No52_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => Delay4No52_out);

   Delay4No53_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => Delay4No53_out);

   Delay4No54_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => Delay4No54_out);

   Delay4No55_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => Delay4No55_out);

   Delay4No56_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => Delay4No56_out);

   Delay4No57_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => Delay4No57_out);

   Delay4No58_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => Delay4No58_out);

   Delay4No59_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => Delay4No59_out);

   Delay4No60_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => Delay4No60_out);

   Delay4No61_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => Delay4No61_out);

   Delay4No62_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => Delay4No62_out);

   Delay4No63_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => Delay4No63_out);

   Delay4No64_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => Delay4No64_out);

   Delay4No65_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => Delay4No65_out);

   Delay4No66_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => Delay4No66_out);

   Delay4No67_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => Delay4No67_out);

   Delay4No68_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => Delay4No68_out);

   Delay4No69_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => Delay4No69_out);

   Delay4No70_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => Delay4No70_out);

   Delay4No71_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => Delay4No71_out);

   Delay4No72_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => Delay4No72_out);

   Delay4No73_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => Delay4No73_out);

   Delay4No74_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => Delay4No74_out);

   Delay4No75_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => Delay4No75_out);

   Delay4No76_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => Delay4No76_out);

   Delay4No77_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => Delay4No77_out);

   Delay4No78_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => Delay4No78_out);

   Delay4No79_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => Delay4No79_out);

   Delay4No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => Delay4No80_out);

   Delay4No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => Delay4No81_out);

   Delay4No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => Delay4No82_out);

   Delay4No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => Delay4No83_out);

   Delay4No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => Delay4No84_out);

   Delay4No85_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => Delay4No85_out);

   Delay4No86_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => Delay4No86_out);

   Delay4No87_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => Delay4No87_out);

   Delay4No88_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => Delay4No88_out);

   Delay4No89_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => Delay4No89_out);

   Delay3No215_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => Delay3No215_out);

   Delay3No216_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => Delay3No216_out);

   Delay3No217_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => Delay3No217_out);

   Delay3No218_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => Delay3No218_out);

   Delay3No219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => Delay3No219_out);

   Delay4No90_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => Delay4No90_out);

   Delay4No91_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => Delay4No91_out);

   Delay4No92_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => Delay4No92_out);

   Delay4No93_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => Delay4No93_out);

   Delay4No94_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => Delay4No94_out);

   Delay4No95_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => Delay4No95_out);

   Delay4No96_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => Delay4No96_out);

   Delay4No97_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => Delay4No97_out);

   Delay4No98_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => Delay4No98_out);

   Delay4No99_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => Delay4No99_out);

   Delay3No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => Delay3No220_out);

   Delay3No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => Delay3No221_out);

   Delay3No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => Delay3No222_out);

   Delay3No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => Delay3No223_out);

   Delay3No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => Delay3No224_out);

   Delay8No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => Delay8No50_out);

   Delay8No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => Delay8No51_out);

   Delay8No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => Delay8No52_out);

   Delay8No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => Delay8No53_out);

   Delay8No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => Delay8No54_out);

   Delay3No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => Delay3No230_out);

   Delay3No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => Delay3No231_out);

   Delay3No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => Delay3No232_out);

   Delay3No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => Delay3No233_out);

   Delay3No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => Delay3No234_out);

   Delay3No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => Delay3No235_out);

   Delay3No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => Delay3No236_out);

   Delay3No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => Delay3No237_out);

   Delay3No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => Delay3No238_out);

   Delay3No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => Delay3No239_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_3_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Add84_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add84_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_Add84_4_impl_0_LUT_out);

   MUX_Add84_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add84_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_Add84_4_impl_1_LUT_out);

   MUX_Subtract135_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract135_4_impl_0_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_Subtract135_4_impl_0_LUT_out);

   MUX_Subtract135_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract135_4_impl_1_LUT_wIn_3_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount61_out,
                 Output => MUX_Subtract135_4_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_0_impl_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_1_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_2_impl_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_3_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_4_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_0_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_1_impl_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_2_impl_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_3_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_4_impl_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add5_1_impl_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add5_2_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add6_4_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add15_4_impl_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_0_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_3_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_4_impl_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_0_impl_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_1_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_2_impl_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_3_impl_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_4_impl_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_0_impl_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_1_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_2_impl_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_3_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_4_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_0_impl_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_1_impl_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_2_impl_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_3_impl_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_4_impl_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add19_2_impl_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add19_3_impl_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add115_1_impl_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add116_0_impl_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add116_1_impl_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add116_2_impl_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_0_impl_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_1_impl_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_2_impl_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add117_3_impl_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add29_3_impl_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add36_4_impl_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add126_0_impl_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add126_4_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add37_2_impl_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_1_impl_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_2_impl_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_3_impl_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add38_0_impl_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add38_1_impl_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add38_2_impl_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add38_3_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_0_impl_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_1_impl_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_2_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_3_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_4_impl_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_0_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_1_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_2_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_3_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_4_impl_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_0_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_1_impl_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_2_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_3_impl_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_4_impl_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_0_impl_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_1_impl_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_2_impl_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_3_impl_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_4_impl_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_0_impl_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_1_impl_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_2_impl_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_3_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_4_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_1_impl_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_2_impl_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_3_impl_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_4_impl_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_0_impl_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_1_impl_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_2_impl_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_3_impl_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_4_impl_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_0_impl_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_1_impl_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_2_impl_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_3_impl_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_4_impl_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_2_impl_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_0_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_1_impl_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_2_impl_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_3_impl_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_0_impl_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_1_impl_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_2_impl_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_3_impl_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_4_impl_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_0_impl_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_1_impl_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_2_impl_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_3_impl_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_4_impl_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_0_impl_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_1_impl_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_2_impl_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_3_impl_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_4_impl_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_0_impl_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_1_impl_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_2_impl_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_3_impl_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_4_impl_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_1_impl_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_2_impl_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_3_impl_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_4_impl_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract5_4_impl_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_0_impl_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_1_impl_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_2_impl_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract6_3_impl_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_0_impl_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_1_impl_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_2_impl_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_3_impl_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product9_4_impl_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_0_impl_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_1_impl_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_2_impl_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_3_impl_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_4_impl_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_0_impl_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_1_impl_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_2_impl_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_3_impl_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract7_4_impl_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_0_impl_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_1_impl_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_2_impl_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_3_impl_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_4_impl_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_0_impl_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_1_impl_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_2_impl_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_3_impl_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_4_impl_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_4_impl_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add50_4_impl_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_0_impl_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_1_impl_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_2_impl_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_3_impl_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product18_4_impl_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_0_impl_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_1_impl_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_2_impl_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_3_impl_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product19_4_impl_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_0_impl_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_1_impl_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_2_impl_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_3_impl_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product28_4_impl_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_0_impl_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_1_impl_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_2_impl_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_3_impl_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product38_4_impl_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_3_impl_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add52_0_impl_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add52_1_impl_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add52_2_impl_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add52_3_impl_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add54_0_impl_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add54_3_impl_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add54_4_impl_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_0_impl_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_1_impl_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_2_impl_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_3_impl_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_4_impl_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_0_impl_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_1_impl_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_2_impl_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_3_impl_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_4_impl_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_0_impl_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_1_impl_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_2_impl_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_3_impl_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_4_impl_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_0_impl_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_1_impl_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_2_impl_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_3_impl_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_4_impl_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract14_4_impl_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract17_0_impl_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract17_1_impl_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_0_impl_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_1_impl_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract18_2_impl_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract19_3_impl_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_0_impl_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_1_impl_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_2_impl_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_4_impl_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract21_0_impl_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract21_1_impl_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract21_2_impl_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract21_3_impl_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract21_4_impl_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add63_4_impl_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_0_impl_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_1_impl_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_2_impl_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_3_impl_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product50_4_impl_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_0_impl_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_1_impl_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_2_impl_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_3_impl_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_4_impl_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_0_impl_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_1_impl_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_2_impl_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_3_impl_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_4_impl_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_0_impl_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_1_impl_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_2_impl_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_3_impl_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_4_impl_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract23_2_impl_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_0_impl_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_1_impl_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_2_impl_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_3_impl_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product124_4_impl_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_0_impl_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_1_impl_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_2_impl_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_3_impl_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_4_impl_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_0_impl_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_1_impl_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_2_impl_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_3_impl_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_4_impl_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_0_impl_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_1_impl_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_2_impl_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_3_impl_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_4_impl_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_0_impl_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_1_impl_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_2_impl_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_3_impl_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_4_impl_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_0_impl_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_1_impl_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_2_impl_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_3_impl_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_4_impl_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_0_impl_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_1_impl_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_2_impl_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_3_impl_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_4_impl_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_0_impl_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_1_impl_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_2_impl_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_3_impl_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_4_impl_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract27_0_impl_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract27_1_impl_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract27_2_impl_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract27_3_impl_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract27_4_impl_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_0_impl_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_1_impl_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_2_impl_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_3_impl_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract42_4_impl_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add84_4_impl_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_0_impl_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_1_impl_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_2_impl_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_3_impl_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract44_4_impl_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract45_3_impl_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_0_impl_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_1_impl_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_2_impl_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_3_impl_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_4_impl_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract47_2_impl_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract47_3_impl_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract47_4_impl_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract52_0_impl_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract52_1_impl_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract52_2_impl_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract52_3_impl_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract52_4_impl_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract112_0_impl_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract112_1_impl_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract112_2_impl_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract112_3_impl_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract112_4_impl_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract56_0_impl_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract56_1_impl_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract56_2_impl_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract56_3_impl_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract60_0_impl_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract60_4_impl_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract126_4_impl_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract135_4_impl_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg930_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg939_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg950_out);
end architecture;

