--------------------------------------------------------------------------------
--                         ModuloCounter_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_4_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of ModuloCounter_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(1 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 3 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid4609136
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid4609136 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid4609136 is
signal XX_m4609137 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m4609137 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m4609137 <= X ;
   YY_m4609137 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid4609140
--                   (IntAdderClassical_33_f500_uid4609142)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid4609140 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid4609140 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid4609136 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid4609140 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid4609136  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f500_uid4609140  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_4_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
         iS_3 when "11",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_3_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_3_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_3_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid4609999_RightShifter
--                (RightShifter_24_by_max_26_F250_uid4610001)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid4609999_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid4609999_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid4610004
--                  (IntAdderAlternative_27_f250_uid4610008)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid4610004 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid4610004 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid4610011
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid4610011 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid4610011 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid4610014
--                   (IntAdderClassical_34_f250_uid4610016)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid4610014 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid4610014 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid4609999
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid4609999 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid4609999 is
   component FPAdd_8_23_uid4609999_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid4610004 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid4610011 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid4610014 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid4609999_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid4610004  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid4610011  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid4610014  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid4609999 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid4609999  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid4612859_RightShifter
--                (RightShifter_24_by_max_26_F250_uid4612861)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid4612859_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid4612859_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid4612864
--                  (IntAdderAlternative_27_f250_uid4612868)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid4612864 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid4612864 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid4612871
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid4612871 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid4612871 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid4612874
--                   (IntAdderClassical_34_f250_uid4612876)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid4612874 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid4612874 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid4612859
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid4612859 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid4612859 is
   component FPAdd_8_23_uid4612859_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid4612864 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid4612871 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid4612874 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid4612859_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid4612864  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid4612871  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid4612874  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid4612859 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid4612859  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 107 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      Y <= s106;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 108 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      Y <= s107;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 99 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      Y <= s98;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 102 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      Y <= s101;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 111 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      Y <= s110;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 103 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      Y <= s102;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 105 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      Y <= s104;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 54 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      Y <= s53;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_72_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 72 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_72_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_72_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      Y <= s71;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 59 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      Y <= s58;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 49 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      Y <= s48;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 69 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      Y <= s68;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      Y <= s60;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 91 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      Y <= s90;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 38 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      Y <= s37;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 80 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      Y <= s79;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      Y <= s55;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 39 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      Y <= s38;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 76 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      Y <= s75;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 85 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      Y <= s84;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 37 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      Y <= s36;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "01" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "10" when "01",
      "00" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "10" when "01",
      "00" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "10" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "10" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "01" when "01",
      "00" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_110_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 110 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_110_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_110_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      Y <= s109;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_89_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 89 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_89_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_89_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      Y <= s88;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 92 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      Y <= s91;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 123 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      Y <= s122;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 67 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      Y <= s66;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_0 : in std_logic_vector(31 downto 0);
          R_U_0 : in std_logic_vector(31 downto 0);
          R_V_0 : in std_logic_vector(31 downto 0);
          R_W_0 : in std_logic_vector(31 downto 0);
          Inv_11_0 : out std_logic_vector(31 downto 0);
          Inv_12_0 : out std_logic_vector(31 downto 0);
          Inv_13_0 : out std_logic_vector(31 downto 0);
          Inv_21_0 : out std_logic_vector(31 downto 0);
          Inv_22_0 : out std_logic_vector(31 downto 0);
          Inv_23_0 : out std_logic_vector(31 downto 0);
          Inv_31_0 : out std_logic_vector(31 downto 0);
          Inv_32_0 : out std_logic_vector(31 downto 0);
          Inv_33_0 : out std_logic_vector(31 downto 0);
          Inv_41_0 : out std_logic_vector(31 downto 0);
          Inv_42_0 : out std_logic_vector(31 downto 0);
          Inv_43_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_4_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(1 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_4_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_3_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_72_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component Delay_34_DelayLength_110_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_89_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount41_out : std_logic_vector(1 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_11_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_12_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_13_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_21_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_22_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_23_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_31_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_32_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_33_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_41_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_42_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_43_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add131_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add131_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add131_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add210_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add210_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add210_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add210_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add210_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add210_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add20_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add20_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add21_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add25_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add25_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add25_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add25_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add28_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add28_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add28_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add28_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add28_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add28_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add28_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add28_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add28_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add71_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add71_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add71_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add81_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add81_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add81_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add81_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add81_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add81_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product112_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product112_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product113_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product113_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product102_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product102_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product131_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product131_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product131_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product131_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product131_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product131_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product131_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product131_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product131_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product371_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product371_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product371_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product381_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product381_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product381_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product381_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product381_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product381_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product391_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product391_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product391_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product411_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product411_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product411_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product411_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product411_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product411_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product421_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product421_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product421_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product421_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product421_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product421_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product421_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product421_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product421_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product441_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product441_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product441_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product441_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product461_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product461_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product461_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product461_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product481_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product481_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product481_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product481_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product511_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product511_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product511_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product511_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product511_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product511_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product511_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product511_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product511_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product521_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product521_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product521_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product521_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product521_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product521_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product521_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product521_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product521_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product57_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product57_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product57_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product57_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product59_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product59_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product59_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product59_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product61_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product61_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product61_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product61_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product62_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product62_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product62_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product63_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product63_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product63_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product63_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product64_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product64_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product64_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product64_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product66_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product66_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product66_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product66_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product67_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product67_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product67_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product68_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product68_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product68_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product711_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product711_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product711_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product711_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product711_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product711_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product711_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product711_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product711_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product70_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product70_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product70_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product70_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product71_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product71_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product71_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product71_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product76_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product76_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product76_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product76_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product911_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product911_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product911_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product911_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract1_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract1_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract5_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract5_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add211_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add211_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add211_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add6_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product14_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product14_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product14_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product26_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product26_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product27_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product27_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product27_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product48_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product48_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product48_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product48_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay112No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay113No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay110No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay110No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Inv_11_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_12_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_13_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_21_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_22_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_23_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_31_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_32_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_33_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_41_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_42_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Inv_43_0_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract5_2_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract5_2_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add9_2_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add9_2_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product48_2_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product48_2_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No1_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No3_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No4_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No5_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay100No1_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No1_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay103No2_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No7_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No2_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No6_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No3_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No4_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay115No5_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay110No_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No8_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay110No2_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No10_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No1_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay114No2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No9_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay112No2_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay113No1_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No11_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No12_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay111No3_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No14_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_12_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_13_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_21_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_22_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_23_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_31_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_32_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_33_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_41_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_42_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_43_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No41_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No1_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add101_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add101_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No1_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No13_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No1_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No26_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No20_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No9_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Add131_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Add131_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No21_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No24_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Add131_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Add131_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No22_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No1_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No18_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No1_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No19_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Add16_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Add16_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No2_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Add210_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Add210_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay68No_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No27_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Add210_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Add210_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No1_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No31_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Add20_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Add20_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No2_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Add21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Add21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No30_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Add21_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Add21_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay12No25_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No1_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No1_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Add23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Add23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Add23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Add23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No1_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Add23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Add23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Add25_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Add25_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No3_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Add25_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Add25_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No1_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Add25_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Add25_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No5_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay17No5_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Add28_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Add28_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Add28_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Add28_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No1_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No1_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Add28_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Add28_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No2_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No32_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Add71_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Add71_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No2_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay71No2_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Add81_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Add81_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Add81_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Add81_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No1_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product113_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product113_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No6_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product113_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product113_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No7_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product113_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product113_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No8_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product102_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product102_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product114_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product114_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No54_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product114_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product114_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No55_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product114_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product114_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product131_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product131_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No9_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product131_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product131_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No10_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product131_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product131_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product371_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product371_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product381_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product381_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product381_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product381_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No58_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product391_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product391_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product411_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product411_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No15_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product411_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product411_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product421_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product421_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product421_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product421_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No16_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Product421_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Product421_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Product441_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Product441_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product441_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product441_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Product441_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Product441_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product461_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product461_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No21_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Product461_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Product461_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Product461_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Product461_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Product481_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Product481_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No24_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product481_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product481_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product481_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product481_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product511_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product511_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No60_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product511_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product511_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No13_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No25_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product511_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product511_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Product521_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Product521_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Product521_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Product521_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Product521_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Product521_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No45_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Product57_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Product57_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Product57_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Product57_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product57_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product57_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product59_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product59_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Product59_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Product59_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Product59_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Product59_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Product61_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Product61_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Product61_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Product61_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Product61_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Product61_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product62_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product62_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Product62_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Product62_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Product62_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Product62_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No44_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Product63_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Product63_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Product63_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Product63_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Product63_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Product63_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product64_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product64_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product64_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product64_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Product64_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Product64_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Product66_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Product66_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Product66_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Product66_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Product66_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Product66_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Product67_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Product67_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Product67_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Product67_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Product67_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Product67_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Product68_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Product68_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Product68_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Product68_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Product68_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Product68_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Product711_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Product711_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Product711_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Product711_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Product711_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Product711_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Product70_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Product70_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No18_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Product70_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Product70_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No19_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Product70_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Product70_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Product71_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Product71_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out_to_Product71_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out_to_Product71_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out_to_Product71_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out_to_Product71_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No23_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out_to_Product76_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out_to_Product76_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out_to_Product76_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out_to_Product76_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out_to_Product76_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out_to_Product76_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out_to_Product911_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out_to_Product911_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out_to_Product911_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out_to_Product911_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out_to_Product911_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out_to_Product911_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No3_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No9_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No4_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No1_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No10_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No5_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No7_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out_to_Subtract1_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out_to_Subtract1_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay18No5_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out_to_Subtract11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out_to_Subtract11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No28_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No27_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No21_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No18_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No22_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No19_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No1_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No8_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No8_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No330_out_to_Subtract5_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No331_out_to_Subtract5_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No20_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No11_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No2_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out_to_Add32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out_to_Add32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out_to_Add32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out_to_Add32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay95No2_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No2_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No14_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out_to_Add211_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out_to_Add211_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay37No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay32No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out_to_Add6_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out_to_Add6_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay51No2_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay57No2_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No54_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out_to_Product11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out_to_Product11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No56_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No350_out_to_Product14_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No351_out_to_Product14_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No352_out_to_Product14_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No353_out_to_Product14_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No46_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No354_out_to_Product14_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No355_out_to_Product14_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No65_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No356_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No357_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No63_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No33_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No358_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No359_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No34_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No49_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No360_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No361_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No362_out_to_Product27_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No363_out_to_Product27_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No364_out_to_Product27_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No365_out_to_Product27_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No366_out_to_Product27_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No367_out_to_Product27_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No368_out_to_Product48_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No369_out_to_Product48_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No370_out_to_Product48_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No371_out_to_Product48_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No372_out_to_Product48_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No373_out_to_Product48_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No374_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No375_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount41_instance: ModuloCounter_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount41_out);
Ldiff_UU_del_1_0_IEEE <= Ldiff_UU_del_1_0;
   Ldiff_UU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_0_out,
                 X => Ldiff_UU_del_1_0_IEEE);
Ldiff_UV_del_1_0_IEEE <= Ldiff_UV_del_1_0;
   Ldiff_UV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_0_out,
                 X => Ldiff_UV_del_1_0_IEEE);
Ldiff_UW_del_1_0_IEEE <= Ldiff_UW_del_1_0;
   Ldiff_UW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_0_out,
                 X => Ldiff_UW_del_1_0_IEEE);
Ldiff_VU_del_1_0_IEEE <= Ldiff_VU_del_1_0;
   Ldiff_VU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_0_out,
                 X => Ldiff_VU_del_1_0_IEEE);
Ldiff_VV_del_1_0_IEEE <= Ldiff_VV_del_1_0;
   Ldiff_VV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_0_out,
                 X => Ldiff_VV_del_1_0_IEEE);
Ldiff_VW_del_1_0_IEEE <= Ldiff_VW_del_1_0;
   Ldiff_VW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_0_out,
                 X => Ldiff_VW_del_1_0_IEEE);
Ldiff_WU_del_1_0_IEEE <= Ldiff_WU_del_1_0;
   Ldiff_WU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_0_out,
                 X => Ldiff_WU_del_1_0_IEEE);
Ldiff_WV_del_1_0_IEEE <= Ldiff_WV_del_1_0;
   Ldiff_WV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_0_out,
                 X => Ldiff_WV_del_1_0_IEEE);
Ldiff_WW_del_1_0_IEEE <= Ldiff_WW_del_1_0;
   Ldiff_WW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_0_out,
                 X => Ldiff_WW_del_1_0_IEEE);
R_U_0_IEEE <= R_U_0;
   R_U_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_0_out,
                 X => R_U_0_IEEE);
R_V_0_IEEE <= R_V_0;
   R_V_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_0_out,
                 X => R_V_0_IEEE);
R_W_0_IEEE <= R_W_0;
   R_W_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_0_out,
                 X => R_W_0_IEEE);

Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_0_impl_out,
                 X => Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg77_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg77_out;
   MUX_Product108_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product108_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg100_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg16_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg114_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
   MUX_Product108_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product108_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product108_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_1_impl_out,
                 X => Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg353_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg5_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product108_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product108_1_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_0_out,
                 Y => Delay1No2_out);

SharedReg390_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
Delay111No1_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast <= Delay111No1_out;
SharedReg9_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product108_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay111No1_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product108_1_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product108_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_2_impl_out,
                 X => Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg377_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg377_out;
SharedReg30_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg353_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product108_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg377_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg30_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product108_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg400_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg400_out;
SharedReg388_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg388_out;
SharedReg109_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg109_out;
   MUX_Product108_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg400_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg388_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg109_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product108_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product110_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_0_impl_out,
                 X => Delay1No6_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg5_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product110_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product110_0_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_0_out,
                 Y => Delay1No6_out);

Delay114No3_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast <= Delay114No3_out;
SharedReg9_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product110_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay114No3_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product110_0_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product110_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_1_impl_out,
                 X => Delay1No8_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast);

SharedReg33_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg353_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg216_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg216_out;
SharedReg275_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg275_out;
   MUX_Product110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg216_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg275_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product110_1_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_0_out,
                 Y => Delay1No8_out);

SharedReg25_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
Delay114No4_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast <= Delay114No4_out;
SharedReg391_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay114No4_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product110_1_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product110_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_2_impl_out,
                 X => Delay1No10_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg91_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg91_out;
SharedReg353_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg91_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product110_2_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_0_out,
                 Y => Delay1No10_out);

SharedReg9_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg386_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
Delay114No5_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast <= Delay114No5_out;
   MUX_Product110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay114No5_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product110_2_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product109_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_0_impl_out,
                 X => Delay1No12_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg215_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg215_out;
SharedReg274_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg274_out;
SharedReg35_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg35_out;
   MUX_Product109_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg274_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg35_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product109_0_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_0_impl_0_out,
                 Y => Delay1No12_out);

SharedReg154_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg391_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg25_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
   MUX_Product109_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product109_0_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_0_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product109_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_1_impl_out,
                 X => Delay1No14_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg353_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg170_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg170_out;
SharedReg280_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg280_out;
   MUX_Product109_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg170_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg280_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product109_1_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_1_impl_0_out,
                 Y => Delay1No14_out);

SharedReg390_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
Delay100No1_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast <= Delay100No1_out;
SharedReg391_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product109_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay100No1_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product109_1_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_1_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product109_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_2_impl_out,
                 X => Delay1No16_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast);

SharedReg213_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg213_out;
SharedReg389_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg353_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product109_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product109_2_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_0_out,
                 Y => Delay1No16_out);

SharedReg391_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg157_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg157_out;
   MUX_Product109_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg157_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product109_2_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product111_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_0_impl_out,
                 X => Delay1No18_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg31_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg278_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg278_out;
SharedReg390_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product111_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg278_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_0_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_0_out,
                 Y => Delay1No18_out);

Delay103No_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast <= Delay103No_out;
SharedReg391_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg390_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product111_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay103No_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_0_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product111_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_1_impl_out,
                 X => Delay1No20_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg353_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg33_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg33_out;
SharedReg389_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg33_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_1_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_0_out,
                 Y => Delay1No20_out);

SharedReg390_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
Delay103No1_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast <= Delay103No1_out;
SharedReg391_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay103No1_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_1_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product111_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_2_impl_out,
                 X => Delay1No22_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg34_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg34_out;
SharedReg276_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg276_out;
SharedReg45_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg45_out;
SharedReg353_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg34_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg276_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg45_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_2_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_0_out,
                 Y => Delay1No22_out);

SharedReg391_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg25_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
Delay103No2_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast <= Delay103No2_out;
   MUX_Product111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay103No2_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_2_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_1_out,
                 Y => Delay1No23_out);

Delay1No24_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast <= Delay1No24_out;
Delay1No25_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast <= Delay1No25_out;
   Product210_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_0_impl_out,
                 X => Delay1No24_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No25_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg35_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg35_out;
SharedReg389_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product210_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg35_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_0_impl_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_0_out,
                 Y => Delay1No24_out);

Delay115No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast <= Delay115No_out;
SharedReg391_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product210_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay115No_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_0_impl_1_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_1_out,
                 Y => Delay1No25_out);

Delay1No26_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast <= Delay1No26_out;
Delay1No27_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast <= Delay1No27_out;
   Product210_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_1_impl_out,
                 X => Delay1No26_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No27_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast);

Delay6No7_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast <= Delay6No7_out;
SharedReg353_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg388_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg388_out;
SharedReg389_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product210_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No7_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg388_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_1_impl_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_0_out,
                 Y => Delay1No26_out);

SharedReg169_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
Delay115No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast <= Delay115No1_out;
SharedReg388_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg388_out;
SharedReg389_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product210_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay115No1_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg388_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_1_impl_1_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_1_out,
                 Y => Delay1No27_out);

Delay1No28_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast <= Delay1No28_out;
Delay1No29_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast <= Delay1No29_out;
   Product210_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_2_impl_out,
                 X => Delay1No28_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No29_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast);

SharedReg39_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg282_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg282_out;
SharedReg390_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg353_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product210_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg282_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_2_impl_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_0_out,
                 Y => Delay1No28_out);

SharedReg391_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg390_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
Delay115No2_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast <= Delay115No2_out;
   MUX_Product210_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay115No2_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_2_impl_1_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_1_out,
                 Y => Delay1No29_out);

Delay1No30_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast <= Delay1No30_out;
Delay1No31_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast <= Delay1No31_out;
   Product310_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_0_impl_out,
                 X => Delay1No30_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No31_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg388_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg389_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
Delay6No6_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast <= Delay6No6_out;
   MUX_Product310_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay6No6_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_0_impl_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_0_out,
                 Y => Delay1No30_out);

Delay115No3_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast <= Delay115No3_out;
SharedReg388_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg389_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg105_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product310_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay115No3_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_0_impl_1_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_1_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Product310_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_1_impl_out,
                 X => Delay1No32_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast);

SharedReg44_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg353_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg16_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product310_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_1_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_0_out,
                 Y => Delay1No32_out);

SharedReg2_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg2_out;
Delay115No4_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast <= Delay115No4_out;
SharedReg24_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product310_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay115No4_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_1_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Product310_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_2_impl_out,
                 X => Delay1No34_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast);

SharedReg388_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg389_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg353_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product310_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_2_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_0_out,
                 Y => Delay1No34_out);

SharedReg388_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg389_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
Delay115No5_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast <= Delay115No5_out;
   MUX_Product310_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay115No5_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_2_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Product410_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_0_impl_out,
                 X => Delay1No36_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg16_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg47_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg47_out;
   MUX_Product410_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg47_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product410_0_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_0_impl_0_out,
                 Y => Delay1No36_out);

Delay110No_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast <= Delay110No_out;
SharedReg24_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg2_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg2_out;
   MUX_Product410_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay110No_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product410_0_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_0_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Product410_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_1_impl_out,
                 X => Delay1No38_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast);

SharedReg48_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg353_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg9_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product410_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product410_1_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_1_impl_0_out,
                 Y => Delay1No38_out);

SharedReg17_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg17_out;
SharedReg128_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg128_out;
SharedReg24_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product410_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg17_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg128_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product410_1_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_1_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Product410_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_2_impl_out,
                 X => Delay1No40_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast);

SharedReg16_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
Delay6No8_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast <= Delay6No8_out;
SharedReg353_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product410_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay6No8_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product410_2_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_2_impl_0_out,
                 Y => Delay1No40_out);

SharedReg24_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg351_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
Delay110No2_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast <= Delay110No2_out;
   MUX_Product410_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg351_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay110No2_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product410_2_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_2_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Product510_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_0_impl_out,
                 X => Delay1No42_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg9_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg51_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg51_out;
   MUX_Product510_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg51_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product510_0_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_0_impl_0_out,
                 Y => Delay1No42_out);

Delay114No_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast <= Delay114No_out;
SharedReg24_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg17_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
   MUX_Product510_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay114No_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product510_0_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_0_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Product510_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_1_impl_out,
                 X => Delay1No44_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast);

Delay2No10_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast <= Delay2No10_out;
SharedReg353_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg16_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product510_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No10_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product510_1_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_1_impl_0_out,
                 Y => Delay1No44_out);

SharedReg6_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg6_out;
Delay114No1_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast <= Delay114No1_out;
SharedReg20_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product510_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay114No1_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product510_1_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_1_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Product510_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_2_impl_out,
                 X => Delay1No46_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast);

SharedReg9_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg55_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg353_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product510_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product510_2_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_2_impl_0_out,
                 Y => Delay1No46_out);

SharedReg24_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg2_out;
Delay114No2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast <= Delay114No2_out;
   MUX_Product510_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay114No2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product510_2_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_2_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Product610_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_0_impl_out,
                 X => Delay1No48_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg16_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
Delay2No9_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast <= Delay2No9_out;
   MUX_Product610_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No9_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product610_0_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_0_out,
                 Y => Delay1No48_out);

SharedReg125_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg125_out;
SharedReg20_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg6_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg6_out;
   MUX_Product610_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg125_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product610_0_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Product610_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_1_impl_out,
                 X => Delay1No50_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast);

SharedReg68_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg353_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg59_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg59_out;
SharedReg389_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product610_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg59_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product610_1_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_0_out,
                 Y => Delay1No50_out);

SharedReg11_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg129_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg129_out;
SharedReg391_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product610_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg129_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product610_1_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Product610_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_2_impl_out,
                 X => Delay1No52_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast);

SharedReg16_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg60_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg60_out;
SharedReg353_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product610_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg60_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product610_2_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_0_out,
                 Y => Delay1No52_out);

SharedReg20_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg17_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
Delay112No2_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast <= Delay112No2_out;
   MUX_Product610_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg17_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay112No2_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product610_2_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product710_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_0_impl_out,
                 X => Delay1No54_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg62_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg389_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg71_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg71_out;
   MUX_Product710_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg71_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product710_0_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_0_impl_0_out,
                 Y => Delay1No54_out);

SharedReg126_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg126_out;
SharedReg391_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg11_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg11_out;
   MUX_Product710_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg126_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product710_0_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_0_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Product710_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_1_impl_out,
                 X => Delay1No56_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast);

Delay2No13_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast <= Delay2No13_out;
SharedReg353_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg63_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg63_out;
SharedReg389_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product710_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No13_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg63_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product710_1_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_0_out,
                 Y => Delay1No56_out);

SharedReg25_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
Delay113No1_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast <= Delay113No1_out;
SharedReg391_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product710_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay113No1_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product710_1_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product710_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_2_impl_out,
                 X => Delay1No58_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast);

SharedReg64_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg64_out;
SharedReg389_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
Delay2No11_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast <= Delay2No11_out;
SharedReg353_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product710_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg64_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No11_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product710_2_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_2_impl_0_out,
                 Y => Delay1No58_out);

SharedReg391_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg6_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg119_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg119_out;
   MUX_Product710_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg6_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg119_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product710_2_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_2_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product810_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_0_impl_out,
                 X => Delay1No60_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg66_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg389_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
Delay2No12_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast <= Delay2No12_out;
   MUX_Product810_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No12_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product810_0_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_0_out,
                 Y => Delay1No60_out);

Delay111No3_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast <= Delay111No3_out;
SharedReg391_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg25_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
   MUX_Product810_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay111No3_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product810_0_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product810_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_1_impl_out,
                 X => Delay1No62_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg353_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg67_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg389_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product810_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg67_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product810_1_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_0_out,
                 Y => Delay1No62_out);

SharedReg17_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg17_out;
SharedReg116_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg116_out;
SharedReg391_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product810_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg17_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg116_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product810_1_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product810_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_2_impl_out,
                 X => Delay1No64_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast);

SharedReg69_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg389_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg83_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg83_out;
SharedReg353_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product810_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg83_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product810_2_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_0_out,
                 Y => Delay1No64_out);

SharedReg391_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg11_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg118_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg118_out;
   MUX_Product810_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg11_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg118_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product810_2_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product910_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_0_impl_out,
                 X => Delay1No66_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast);

SharedReg353_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg70_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg70_out;
SharedReg389_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg86_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg86_out;
   MUX_Product910_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg70_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg86_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product910_0_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_0_impl_0_out,
                 Y => Delay1No66_out);

SharedReg142_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg391_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg17_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg17_out;
   MUX_Product910_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg17_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product910_0_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_0_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product910_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_1_impl_out,
                 X => Delay1No68_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg353_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg353_out;
SharedReg5_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product910_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg353_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product910_1_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_0_out,
                 Y => Delay1No68_out);

SharedReg21_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg145_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg145_out;
SharedReg20_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product910_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product910_1_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product910_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_2_impl_out,
                 X => Delay1No70_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast);

SharedReg75_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg389_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
Delay2No14_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast <= Delay2No14_out;
SharedReg353_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg353_out;
   MUX_Product910_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No14_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg353_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product910_2_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_2_impl_0_out,
                 Y => Delay1No70_out);

SharedReg391_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg25_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg139_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg139_out;
   MUX_Product910_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg139_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product910_2_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_2_impl_1_out,
                 Y => Delay1No71_out);
   Inv_11_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_0_IEEE,
                 X => Delay1No72_out);
Inv_11_0 <= Inv_11_0_IEEE;

SharedReg31_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast <= SharedReg31_out;
SharedReg33_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg34_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast <= SharedReg34_out;
   MUX_Inv_11_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg31_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg34_out_to_MUX_Inv_11_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_11_0_0_LUT_out,
                 oMux => MUX_Inv_11_0_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_11_0_0_out,
                 Y => Delay1No72_out);
   Inv_12_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_0_IEEE,
                 X => Delay1No73_out);
Inv_12_0 <= Inv_12_0_IEEE;

SharedReg35_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg36_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast <= SharedReg36_out;
SharedReg39_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast <= SharedReg39_out;
   MUX_Inv_12_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg39_out_to_MUX_Inv_12_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_12_0_0_LUT_out,
                 oMux => MUX_Inv_12_0_0_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_12_0_0_out,
                 Y => Delay1No73_out);
   Inv_13_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_0_IEEE,
                 X => Delay1No74_out);
Inv_13_0 <= Inv_13_0_IEEE;

SharedReg51_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast <= SharedReg51_out;
SharedReg52_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast <= SharedReg52_out;
SharedReg55_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast <= SharedReg55_out;
   MUX_Inv_13_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg51_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg52_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_Inv_13_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_13_0_0_LUT_out,
                 oMux => MUX_Inv_13_0_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_13_0_0_out,
                 Y => Delay1No74_out);
   Inv_21_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_0_IEEE,
                 X => Delay1No75_out);
Inv_21_0 <= Inv_21_0_IEEE;

SharedReg56_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg59_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast <= SharedReg59_out;
SharedReg60_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast <= SharedReg60_out;
   MUX_Inv_21_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg59_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg60_out_to_MUX_Inv_21_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_21_0_0_LUT_out,
                 oMux => MUX_Inv_21_0_0_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_21_0_0_out,
                 Y => Delay1No75_out);
   Inv_22_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_0_IEEE,
                 X => Delay1No76_out);
Inv_22_0 <= Inv_22_0_IEEE;

SharedReg62_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast <= SharedReg62_out;
SharedReg63_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast <= SharedReg63_out;
SharedReg64_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast <= SharedReg64_out;
   MUX_Inv_22_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg62_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg63_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg64_out_to_MUX_Inv_22_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_22_0_0_LUT_out,
                 oMux => MUX_Inv_22_0_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_22_0_0_out,
                 Y => Delay1No76_out);
   Inv_23_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_0_IEEE,
                 X => Delay1No77_out);
Inv_23_0 <= Inv_23_0_IEEE;

SharedReg66_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg67_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast <= SharedReg67_out;
SharedReg69_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast <= SharedReg69_out;
   MUX_Inv_23_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg67_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg69_out_to_MUX_Inv_23_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_23_0_0_LUT_out,
                 oMux => MUX_Inv_23_0_0_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_23_0_0_out,
                 Y => Delay1No77_out);
   Inv_31_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_0_IEEE,
                 X => Delay1No78_out);
Inv_31_0 <= Inv_31_0_IEEE;

SharedReg70_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg72_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg75_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast <= SharedReg75_out;
   MUX_Inv_31_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg75_out_to_MUX_Inv_31_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_31_0_0_LUT_out,
                 oMux => MUX_Inv_31_0_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_31_0_0_out,
                 Y => Delay1No78_out);
   Inv_32_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_0_IEEE,
                 X => Delay1No79_out);
Inv_32_0 <= Inv_32_0_IEEE;

SharedReg76_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast <= SharedReg76_out;
SharedReg79_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast <= SharedReg79_out;
SharedReg82_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast <= SharedReg82_out;
   MUX_Inv_32_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg76_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg79_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg82_out_to_MUX_Inv_32_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_32_0_0_LUT_out,
                 oMux => MUX_Inv_32_0_0_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_32_0_0_out,
                 Y => Delay1No79_out);
   Inv_33_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_0_IEEE,
                 X => Delay1No80_out);
Inv_33_0 <= Inv_33_0_IEEE;

SharedReg85_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast <= SharedReg85_out;
SharedReg88_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast <= SharedReg88_out;
SharedReg90_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
   MUX_Inv_33_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg85_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg88_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg90_out_to_MUX_Inv_33_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_33_0_0_LUT_out,
                 oMux => MUX_Inv_33_0_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_33_0_0_out,
                 Y => Delay1No80_out);
   Inv_41_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_0_IEEE,
                 X => Delay1No81_out);
Inv_41_0 <= Inv_41_0_IEEE;

SharedReg93_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast <= SharedReg93_out;
SharedReg95_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg96_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast <= SharedReg96_out;
   MUX_Inv_41_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg93_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg96_out_to_MUX_Inv_41_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_41_0_0_LUT_out,
                 oMux => MUX_Inv_41_0_0_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_41_0_0_out,
                 Y => Delay1No81_out);
   Inv_42_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_0_IEEE,
                 X => Delay1No82_out);
Inv_42_0 <= Inv_42_0_IEEE;

SharedReg41_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg44_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast <= SharedReg44_out;
SharedReg45_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast <= SharedReg45_out;
   MUX_Inv_42_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg44_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg45_out_to_MUX_Inv_42_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_42_0_0_LUT_out,
                 oMux => MUX_Inv_42_0_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_42_0_0_out,
                 Y => Delay1No82_out);
   Inv_43_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_0_IEEE,
                 X => Delay1No83_out);
Inv_43_0 <= Inv_43_0_IEEE;

SharedReg47_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast <= SharedReg47_out;
SharedReg48_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast <= SharedReg48_out;
SharedReg49_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast <= SharedReg49_out;
   MUX_Inv_43_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg48_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg49_out_to_MUX_Inv_43_0_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Inv_43_0_0_LUT_out,
                 oMux => MUX_Inv_43_0_0_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Inv_43_0_0_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_0_impl_out,
                 X => Delay1No84_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast);

SharedReg230_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg230_out;
Delay14No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast <= Delay14No_out;
SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg221_out;
SharedReg243_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
   MUX_Add30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay14No_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg221_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add30_0_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_0_out,
                 Y => Delay1No84_out);

SharedReg215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg332_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg332_out;
SharedReg338_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg304_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg304_out;
   MUX_Add30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg332_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg338_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg304_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add30_0_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_1_impl_out,
                 X => Delay1No86_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg245_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg245_out;
SharedReg232_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg232_out;
Delay17No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast <= Delay17No1_out;
SharedReg44_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg44_out;
   MUX_Add30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg245_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg232_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay17No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add30_1_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_0_out,
                 Y => Delay1No86_out);

SharedReg306_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg306_out;
SharedReg224_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg224_out;
SharedReg132_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg132_out;
SharedReg127_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg127_out;
   MUX_Add30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg306_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg224_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg132_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg127_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add30_1_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add30_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_2_impl_out,
                 X => Delay1No88_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast);

Delay36No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast <= Delay36No1_out;
Delay32No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast <= Delay32No1_out;
SharedReg246_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg246_out;
SharedReg233_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg233_out;
   MUX_Add30_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay36No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay32No1_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg246_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg233_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add30_2_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_0_out,
                 Y => Delay1No88_out);

SharedReg159_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg159_out;
SharedReg110_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg110_out;
SharedReg307_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg307_out;
Delay2No41_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast <= Delay2No41_out;
   MUX_Add30_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg159_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg307_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No41_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add30_2_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add110_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_1_impl_out,
                 X => Delay1No90_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast);

Delay32No_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast <= Delay32No_out;
SharedReg15_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg176_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg176_out;
Delay36No_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast <= Delay36No_out;
   MUX_Add110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay32No_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg176_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay36No_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add110_1_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_1_impl_0_out,
                 Y => Delay1No90_out);

SharedReg342_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg342_out;
SharedReg381_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg381_out;
SharedReg333_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg333_out;
SharedReg167_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg167_out;
   MUX_Add110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg342_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg381_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg333_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg167_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add110_1_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_1_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add110_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_2_impl_out,
                 X => Delay1No92_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast);

Delay14No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast <= Delay14No2_out;
Delay51No1_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast <= Delay51No1_out;
SharedReg276_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg276_out;
SharedReg254_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg254_out;
   MUX_Add110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay14No2_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay51No1_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg276_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg254_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add110_2_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_0_out,
                 Y => Delay1No92_out);

SharedReg334_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg334_out;
SharedReg334_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg334_out;
SharedReg282_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg282_out;
SharedReg335_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg335_out;
   MUX_Add110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg334_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg334_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg282_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg335_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add110_2_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add101_2_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add101_2_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add101_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_2_impl_out,
                 X => Delay1No94_out_to_Add101_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add101_2_impl_parent_implementedSystem_port_1_cast);

Delay27No1_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_1_cast <= Delay27No1_out;
SharedReg34_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg34_out;
SharedReg27_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg234_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg234_out;
   MUX_Add101_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay27No1_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg34_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg27_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg234_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add101_2_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_2_impl_0_out,
                 Y => Delay1No94_out);

SharedReg155_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg155_out;
Delay11No13_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_2_cast <= Delay11No13_out;
SharedReg34_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg34_out;
SharedReg213_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg213_out;
   MUX_Add101_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg155_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay11No13_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg34_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg213_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add101_2_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_2_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add111_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_1_impl_out,
                 X => Delay1No96_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast);

Delay51No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast <= Delay51No_out;
SharedReg27_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg27_out;
Delay15No1_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast <= Delay15No1_out;
SharedReg225_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg225_out;
   MUX_Add111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay51No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay15No1_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg225_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add111_1_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_0_out,
                 Y => Delay1No96_out);

SharedReg338_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg338_out;
SharedReg170_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg170_out;
SharedReg334_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg334_out;
SharedReg339_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg339_out;
   MUX_Add111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg338_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg170_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg334_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg339_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add111_1_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add111_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_2_impl_out,
                 X => Delay1No98_out_to_Add111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg303_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg303_out;
SharedReg228_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg228_out;
Delay8No26_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_3_cast <= Delay8No26_out;
SharedReg252_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg252_out;
   MUX_Add111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg303_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg228_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay8No26_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Add111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add111_2_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_2_impl_0_out,
                 Y => Delay1No98_out);

SharedReg341_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg341_out;
SharedReg341_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg341_out;
SharedReg340_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg340_out;
Delay12No20_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_4_cast <= Delay12No20_out;
   MUX_Add111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg341_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg340_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay12No20_out_to_MUX_Add111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add111_2_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_2_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add121_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_0_impl_out,
                 X => Delay1No100_out_to_Add121_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add121_0_impl_parent_implementedSystem_port_1_cast);

SharedReg235_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg235_out;
Delay15No_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast <= Delay15No_out;
SharedReg47_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg47_out;
SharedReg274_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg274_out;
   MUX_Add121_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg235_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg47_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg274_out_to_MUX_Add121_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add121_0_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_0_impl_0_out,
                 Y => Delay1No100_out);

SharedReg256_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg333_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg333_out;
Delay5No9_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast <= Delay5No9_out;
SharedReg278_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg278_out;
   MUX_Add121_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay5No9_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg278_out_to_MUX_Add121_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add121_0_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_0_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add121_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_1_impl_out,
                 X => Delay1No102_out_to_Add121_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add121_1_impl_parent_implementedSystem_port_1_cast);

SharedReg275_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg275_out;
SharedReg245_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg245_out;
SharedReg196_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg196_out;
SharedReg328_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg328_out;
   MUX_Add121_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg275_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg245_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg196_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg328_out_to_MUX_Add121_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add121_1_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_1_impl_0_out,
                 Y => Delay1No102_out);

SharedReg280_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg280_out;
SharedReg258_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg258_out;
SharedReg205_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg205_out;
SharedReg333_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg333_out;
   MUX_Add121_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg280_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg258_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg205_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg333_out_to_MUX_Add121_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add121_1_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_1_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Add131_0_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Add131_0_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Add131_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add131_0_impl_out,
                 X => Delay1No104_out_to_Add131_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Add131_0_impl_parent_implementedSystem_port_1_cast);

Delay10No21_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_1_cast <= Delay10No21_out;
Delay17No_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_2_cast <= Delay17No_out;
SharedReg325_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg325_out;
Delay8No24_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_4_cast <= Delay8No24_out;
   MUX_Add131_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay10No21_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay17No_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg325_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay8No24_out_to_MUX_Add131_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add131_0_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_0_impl_0_out,
                 Y => Delay1No104_out);

SharedReg337_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg337_out;
SharedReg130_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg332_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg332_out;
SharedReg337_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg337_out;
   MUX_Add131_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg337_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg332_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg337_out_to_MUX_Add131_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add131_0_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_0_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Add131_1_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Add131_1_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Add131_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add131_1_impl_out,
                 X => Delay1No106_out_to_Add131_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Add131_1_impl_parent_implementedSystem_port_1_cast);

SharedReg251_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg251_out;
Delay10No22_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_2_cast <= Delay10No22_out;
SharedReg44_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg44_out;
Delay16No1_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_4_cast <= Delay16No1_out;
   MUX_Add131_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg251_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay10No22_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg44_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay16No1_out_to_MUX_Add131_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add131_1_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_1_impl_0_out,
                 Y => Delay1No106_out);

SharedReg336_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg336_out;
SharedReg339_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg339_out;
SharedReg48_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg48_out;
SharedReg336_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg336_out;
   MUX_Add131_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg336_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg339_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg48_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg336_out_to_MUX_Add131_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add131_1_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add131_1_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Add16_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_0_impl_out,
                 X => Delay1No108_out_to_Add16_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Add16_0_impl_parent_implementedSystem_port_1_cast);

SharedReg255_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg255_out;
SharedReg203_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg203_out;
Delay16No_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast <= Delay16No_out;
SharedReg308_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg308_out;
   MUX_Add16_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg255_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg203_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay16No_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg308_out_to_MUX_Add16_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_0_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_0_impl_0_out,
                 Y => Delay1No108_out);

Delay12No18_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast <= Delay12No18_out;
SharedReg210_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg210_out;
SharedReg337_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg337_out;
SharedReg314_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg314_out;
   MUX_Add16_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No18_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg210_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg337_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg314_out_to_MUX_Add16_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_0_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_0_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Add16_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_1_impl_out,
                 X => Delay1No110_out_to_Add16_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Add16_1_impl_parent_implementedSystem_port_1_cast);

SharedReg309_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg309_out;
SharedReg261_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg261_out;
SharedReg184_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg184_out;
Delay68No1_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast <= Delay68No1_out;
   MUX_Add16_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg309_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg261_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg184_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay68No1_out_to_MUX_Add16_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_1_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_1_impl_0_out,
                 Y => Delay1No110_out);

SharedReg316_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg316_out;
Delay12No19_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast <= Delay12No19_out;
SharedReg159_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg159_out;
SharedReg161_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg161_out;
   MUX_Add16_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg316_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay12No19_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg159_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg161_out_to_MUX_Add16_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_1_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_1_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Add16_2_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Add16_2_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Add16_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_2_impl_out,
                 X => Delay1No112_out_to_Add16_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Add16_2_impl_parent_implementedSystem_port_1_cast);

Delay17No2_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_1_cast <= Delay17No2_out;
SharedReg55_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg55_out;
SharedReg311_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg311_out;
SharedReg198_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg198_out;
   MUX_Add16_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay17No2_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg311_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg198_out_to_MUX_Add16_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_2_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_2_impl_0_out,
                 Y => Delay1No112_out);

SharedReg117_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg152_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg317_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg50_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg50_out;
   MUX_Add16_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg317_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg50_out_to_MUX_Add16_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_2_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_2_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Add210_0_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Add210_0_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Add210_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add210_0_impl_out,
                 X => Delay1No114_out_to_Add210_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Add210_0_impl_parent_implementedSystem_port_1_cast);

SharedReg193_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg193_out;
SharedReg47_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg47_out;
Delay68No_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_3_cast <= Delay68No_out;
SharedReg222_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg222_out;
   MUX_Add210_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg193_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg47_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay68No_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg222_out_to_MUX_Add210_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add210_0_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add210_0_impl_0_out,
                 Y => Delay1No114_out);

SharedReg42_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg51_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg51_out;
Delay3No27_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_3_cast <= Delay3No27_out;
SharedReg338_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg338_out;
   MUX_Add210_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg51_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No27_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg338_out_to_MUX_Add210_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add210_0_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add210_0_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Add210_1_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Add210_1_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Add210_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add210_1_impl_out,
                 X => Delay1No116_out_to_Add210_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Add210_1_impl_parent_implementedSystem_port_1_cast);

SharedReg226_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg226_out;
SharedReg196_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg196_out;
Delay11No1_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_3_cast <= Delay11No1_out;
Delay90No1_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_4_cast <= Delay90No1_out;
   MUX_Add210_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg196_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay11No1_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay90No1_out_to_MUX_Add210_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add210_1_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add210_1_impl_0_out,
                 Y => Delay1No116_out);

SharedReg339_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg339_out;
SharedReg37_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg336_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg336_out;
Delay3No31_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_4_cast <= Delay3No31_out;
   MUX_Add210_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg339_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg336_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No31_out_to_MUX_Add210_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add210_1_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add210_1_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Add20_2_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Add20_2_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Add20_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add20_2_impl_out,
                 X => Delay1No118_out_to_Add20_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Add20_2_impl_parent_implementedSystem_port_1_cast);

SharedReg201_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg201_out;
SharedReg330_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg330_out;
Delay18No2_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_3_cast <= Delay18No2_out;
SharedReg220_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg220_out;
   MUX_Add20_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg201_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg330_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay18No2_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg220_out_to_MUX_Add20_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add20_2_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_2_impl_0_out,
                 Y => Delay1No118_out);

SharedReg207_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg207_out;
SharedReg335_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg335_out;
SharedReg341_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg341_out;
SharedReg137_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg137_out;
   MUX_Add20_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg207_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg335_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg341_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg137_out_to_MUX_Add20_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add20_2_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add20_2_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Add21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Add21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Add21_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add21_0_impl_out,
                 X => Delay1No120_out_to_Add21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Add21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg223_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg223_out;
SharedReg181_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg181_out;
Delay90No_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_3_cast <= Delay90No_out;
SharedReg279_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg279_out;
   MUX_Add21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg223_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg181_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay90No_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg279_out_to_MUX_Add21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add21_0_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_0_impl_0_out,
                 Y => Delay1No120_out);

SharedReg134_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg158_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg158_out;
Delay3No30_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_3_cast <= Delay3No30_out;
SharedReg332_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg332_out;
   MUX_Add21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg158_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No30_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg332_out_to_MUX_Add21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add21_0_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_0_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Add21_1_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Add21_1_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Add21_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add21_1_impl_out,
                 X => Delay1No122_out_to_Add21_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Add21_1_impl_parent_implementedSystem_port_1_cast);

Delay12No25_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_1_cast <= Delay12No25_out;
Delay21No1_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_2_cast <= Delay21No1_out;
SharedReg74_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
Delay87No1_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_4_cast <= Delay87No1_out;
   MUX_Add21_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay12No25_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay21No1_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg74_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay87No1_out_to_MUX_Add21_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add21_1_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_1_impl_0_out,
                 Y => Delay1No122_out);

SharedReg333_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg333_out;
SharedReg135_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg135_out;
SharedReg339_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg339_out;
SharedReg136_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg136_out;
   MUX_Add21_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg333_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg135_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg339_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg136_out_to_MUX_Add21_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add21_1_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_1_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Add23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Add23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Add23_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_0_impl_out,
                 X => Delay1No124_out_to_Add23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Add23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg283_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg283_out;
Delay11No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_2_cast <= Delay11No_out;
Delay87No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_3_cast <= Delay87No_out;
SharedReg62_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg62_out;
   MUX_Add23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg283_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay11No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay87No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add23_0_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_0_impl_0_out,
                 Y => Delay1No124_out);

SharedReg131_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg337_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg337_out;
SharedReg141_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg141_out;
SharedReg66_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg66_out;
   MUX_Add23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg337_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg141_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg66_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add23_0_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_0_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Add23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Add23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Add23_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_1_impl_out,
                 X => Delay1No126_out_to_Add23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Add23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg59_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg59_out;
SharedReg288_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg288_out;
SharedReg368_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg368_out;
Delay95No1_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_4_cast <= Delay95No1_out;
   MUX_Add23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg59_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg288_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg368_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay95No1_out_to_MUX_Add23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add23_1_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_1_impl_0_out,
                 Y => Delay1No126_out);

SharedReg63_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg123_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg123_out;
SharedReg110_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg110_out;
SharedReg144_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg144_out;
   MUX_Add23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg110_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg144_out_to_MUX_Add23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add23_1_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_1_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Add23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Add23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Add23_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_2_impl_out,
                 X => Delay1No128_out_to_Add23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Add23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg49_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg200_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg200_out;
SharedReg277_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg277_out;
SharedReg282_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg282_out;
   MUX_Add23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg200_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg277_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg282_out_to_MUX_Add23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add23_2_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_2_impl_0_out,
                 Y => Delay1No128_out);

SharedReg55_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg55_out;
SharedReg340_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg340_out;
SharedReg335_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg335_out;
SharedReg138_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg138_out;
   MUX_Add23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg55_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg340_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg335_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg138_out_to_MUX_Add23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add23_2_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_2_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Add25_0_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Add25_0_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Add25_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add25_0_impl_out,
                 X => Delay1No130_out_to_Add25_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Add25_0_impl_parent_implementedSystem_port_1_cast);

Delay17No3_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_1_cast <= Delay17No3_out;
SharedReg78_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg78_out;
Delay95No_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_3_cast <= Delay95No_out;
SharedReg93_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg93_out;
   MUX_Add25_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay17No3_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay95No_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg93_out_to_MUX_Add25_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add25_0_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_0_impl_0_out,
                 Y => Delay1No130_out);

SharedReg140_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg140_out;
SharedReg338_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg148_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg148_out;
SharedReg187_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg187_out;
   MUX_Add25_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg140_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg148_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg187_out_to_MUX_Add25_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add25_0_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_0_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Add25_1_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Add25_1_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Add25_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add25_1_impl_out,
                 X => Delay1No132_out_to_Add25_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Add25_1_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg281_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg281_out;
Delay37No1_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_3_cast <= Delay37No1_out;
SharedReg362_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg362_out;
   MUX_Add25_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg281_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay37No1_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg362_out_to_MUX_Add25_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add25_1_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_1_impl_0_out,
                 Y => Delay1No132_out);

SharedReg95_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg143_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg143_out;
SharedReg102_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg102_out;
SharedReg149_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg149_out;
   MUX_Add25_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg143_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg102_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg149_out_to_MUX_Add25_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add25_1_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_1_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Add25_2_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Add25_2_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Add25_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add25_2_impl_out,
                 X => Delay1No134_out_to_Add25_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Add25_2_impl_parent_implementedSystem_port_1_cast);

Delay14No5_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_1_cast <= Delay14No5_out;
SharedReg364_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg364_out;
SharedReg69_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg69_out;
Delay17No5_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_4_cast <= Delay17No5_out;
   MUX_Add25_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay14No5_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg364_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg69_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay17No5_out_to_MUX_Add25_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add25_2_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_2_impl_0_out,
                 Y => Delay1No134_out);

SharedReg162_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg162_out;
SharedReg165_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg75_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg75_out;
SharedReg150_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg150_out;
   MUX_Add25_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg162_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg75_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg150_out_to_MUX_Add25_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add25_2_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add25_2_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Add28_0_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Add28_0_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Add28_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add28_0_impl_out,
                 X => Delay1No136_out_to_Add28_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Add28_0_impl_parent_implementedSystem_port_1_cast);

Delay20No_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_1_cast <= Delay20No_out;
SharedReg360_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg360_out;
SharedReg355_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg355_out;
Delay71No_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_4_cast <= Delay71No_out;
   MUX_Add28_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay20No_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg360_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg355_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay71No_out_to_MUX_Add28_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add28_0_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add28_0_impl_0_out,
                 Y => Delay1No136_out);

SharedReg332_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg332_out;
SharedReg342_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg342_out;
SharedReg158_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg158_out;
SharedReg342_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg342_out;
   MUX_Add28_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg332_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg342_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg158_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg342_out_to_MUX_Add28_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add28_0_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add28_0_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Add28_1_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Add28_1_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Add28_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add28_1_impl_out,
                 X => Delay1No138_out_to_Add28_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Add28_1_impl_parent_implementedSystem_port_1_cast);

Delay71No1_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_1_cast <= Delay71No1_out;
Delay20No1_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_2_cast <= Delay20No1_out;
SharedReg_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg_out;
SharedReg369_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg369_out;
   MUX_Add28_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay71No1_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay20No1_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg369_out_to_MUX_Add28_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add28_1_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add28_1_impl_0_out,
                 Y => Delay1No138_out);

SharedReg168_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg168_out;
SharedReg336_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg336_out;
SharedReg377_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg377_out;
SharedReg155_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg155_out;
   MUX_Add28_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg168_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg336_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg377_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg155_out_to_MUX_Add28_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add28_1_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add28_1_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Add28_2_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Add28_2_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Add28_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add28_2_impl_out,
                 X => Delay1No140_out_to_Add28_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Add28_2_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
Delay90No2_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_2_cast <= Delay90No2_out;
SharedReg191_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg191_out;
Delay20No2_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_4_cast <= Delay20No2_out;
   MUX_Add28_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay90No2_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg191_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay20No2_out_to_MUX_Add28_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add28_2_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add28_2_impl_0_out,
                 Y => Delay1No140_out);

SharedReg335_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg335_out;
Delay3No32_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_2_cast <= Delay3No32_out;
SharedReg177_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg177_out;
SharedReg334_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg334_out;
   MUX_Add28_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg335_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No32_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg177_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg334_out_to_MUX_Add28_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add28_2_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add28_2_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Add71_2_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Add71_2_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Add71_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add71_2_impl_out,
                 X => Delay1No142_out_to_Add71_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Add71_2_impl_parent_implementedSystem_port_1_cast);

SharedReg92_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
Delay87No2_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_2_cast <= Delay87No2_out;
Delay71No2_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_3_cast <= Delay71No2_out;
SharedReg201_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg201_out;
   MUX_Add71_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay87No2_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay71No2_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg201_out_to_MUX_Add71_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add71_2_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add71_2_impl_0_out,
                 Y => Delay1No142_out);

SharedReg340_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg163_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg163_out;
SharedReg350_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg350_out;
SharedReg208_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg208_out;
   MUX_Add71_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg163_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg350_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg208_out_to_MUX_Add71_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add71_2_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add71_2_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Add81_0_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Add81_0_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Add81_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add81_0_impl_out,
                 X => Delay1No144_out_to_Add81_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Add81_0_impl_parent_implementedSystem_port_1_cast);

SharedReg203_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg203_out;
Delay37No_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_2_cast <= Delay37No_out;
SharedReg366_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg366_out;
Delay73No_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_4_cast <= Delay73No_out;
   MUX_Add81_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg203_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay37No_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg366_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay73No_out_to_MUX_Add81_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add81_0_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add81_0_impl_0_out,
                 Y => Delay1No144_out);

SharedReg204_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg204_out;
SharedReg104_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg104_out;
SharedReg167_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg167_out;
SharedReg134_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg134_out;
   MUX_Add81_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg204_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg167_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg134_out_to_MUX_Add81_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add81_0_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add81_0_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Add81_1_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Add81_1_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Add81_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add81_1_impl_out,
                 X => Delay1No146_out_to_Add81_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Add81_1_impl_parent_implementedSystem_port_1_cast);

Delay73No1_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_1_cast <= Delay73No1_out;
SharedReg205_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg15_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg15_out;
SharedReg310_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg310_out;
   MUX_Add81_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay73No1_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg15_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg310_out_to_MUX_Add81_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add81_1_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add81_1_impl_0_out,
                 Y => Delay1No146_out);

SharedReg132_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg197_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg197_out;
SharedReg382_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg382_out;
SharedReg107_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg107_out;
   MUX_Add81_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg197_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg382_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg107_out_to_MUX_Add81_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add81_1_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add81_1_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product112_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product112_1_impl_out,
                 X => Delay1No148_out_to_Product112_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product112_1_impl_parent_implementedSystem_port_1_cast);

SharedReg73_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg30_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg1_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product112_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product112_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product112_1_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_1_impl_0_out,
                 Y => Delay1No148_out);

SharedReg111_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg388_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg16_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product112_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product112_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product112_1_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product112_1_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product113_0_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product113_0_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product113_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_0_impl_out,
                 X => Delay1No150_out_to_Product113_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product113_0_impl_parent_implementedSystem_port_1_cast);

Delay3No6_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No6_out;
SharedReg1_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product113_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No6_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product113_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product113_0_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_0_impl_0_out,
                 Y => Delay1No150_out);

SharedReg18_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg20_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product113_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product113_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product113_0_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_0_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product113_1_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product113_1_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product113_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_1_impl_out,
                 X => Delay1No152_out_to_Product113_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product113_1_impl_parent_implementedSystem_port_1_cast);

SharedReg54_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg54_out;
Delay3No7_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_2_cast <= Delay3No7_out;
SharedReg5_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product113_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No7_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product113_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product113_1_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_1_impl_0_out,
                 Y => Delay1No152_out);

SharedReg6_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg18_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product113_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product113_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product113_1_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_1_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product113_2_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product113_2_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product113_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product113_2_impl_out,
                 X => Delay1No154_out_to_Product113_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product113_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg192_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg192_out;
Delay3No8_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_4_cast <= Delay3No8_out;
   MUX_Product113_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg192_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No8_out_to_MUX_Product113_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product113_2_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_2_impl_0_out,
                 Y => Delay1No154_out);

SharedReg20_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg21_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg18_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg18_out;
   MUX_Product113_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg21_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg18_out_to_MUX_Product113_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product113_2_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product113_2_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product102_0_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product102_0_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product102_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_0_impl_out,
                 X => Delay1No156_out_to_Product102_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product102_0_impl_parent_implementedSystem_port_1_cast);

SharedReg287_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg287_out;
SharedReg5_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg58_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg58_out;
   MUX_Product102_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg287_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg58_out_to_MUX_Product102_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product102_0_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_0_impl_0_out,
                 Y => Delay1No156_out);

SharedReg397_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg24_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg6_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg6_out;
   MUX_Product102_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Product102_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product102_0_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_0_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product102_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_1_impl_out,
                 X => Delay1No158_out_to_Product102_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product102_1_impl_parent_implementedSystem_port_1_cast);

SharedReg189_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg294_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg294_out;
SharedReg95_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg389_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product102_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg294_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product102_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product102_1_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_1_impl_0_out,
                 Y => Delay1No158_out);

SharedReg21_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg397_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg391_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product102_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product102_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product102_1_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_1_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product102_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product102_2_impl_out,
                 X => Delay1No160_out_to_Product102_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product102_2_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg286_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg286_out;
   MUX_Product102_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg286_out_to_MUX_Product102_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product102_2_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_2_impl_0_out,
                 Y => Delay1No160_out);

SharedReg24_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg397_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product102_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product102_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product102_2_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product102_2_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product114_0_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product114_0_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product114_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_0_impl_out,
                 X => Delay1No162_out_to_Product114_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product114_0_impl_parent_implementedSystem_port_1_cast);

Delay7No54_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_1_cast <= Delay7No54_out;
SharedReg5_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg94_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg94_out;
   MUX_Product114_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No54_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg94_out_to_MUX_Product114_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_0_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_0_impl_0_out,
                 Y => Delay1No162_out);

SharedReg115_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg20_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg21_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
   MUX_Product114_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Product114_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_0_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_0_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product114_1_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product114_1_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product114_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_1_impl_out,
                 X => Delay1No164_out_to_Product114_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product114_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
Delay7No55_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_2_cast <= Delay7No55_out;
SharedReg1_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product114_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay7No55_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product114_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_1_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_1_impl_0_out,
                 Y => Delay1No164_out);

SharedReg390_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg112_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg20_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product114_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product114_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_1_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_1_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product114_2_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product114_2_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product114_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_2_impl_out,
                 X => Delay1No166_out_to_Product114_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product114_2_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg97_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg97_out;
SharedReg46_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg46_out;
   MUX_Product114_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg97_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg46_out_to_MUX_Product114_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_2_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_2_impl_0_out,
                 Y => Delay1No166_out);

SharedReg20_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg17_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg17_out;
SharedReg387_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
   MUX_Product114_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg17_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg387_out_to_MUX_Product114_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_2_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_2_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product131_0_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product131_0_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product131_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product131_0_impl_out,
                 X => Delay1No168_out_to_Product131_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product131_0_impl_parent_implementedSystem_port_1_cast);

Delay3No9_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No9_out;
SharedReg187_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg187_out;
SharedReg389_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg172_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg172_out;
   MUX_Product131_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No9_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg187_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg172_out_to_MUX_Product131_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product131_0_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product131_0_impl_0_out,
                 Y => Delay1No168_out);

SharedReg7_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg7_out;
SharedReg391_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg21_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
   MUX_Product131_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg7_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Product131_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product131_0_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product131_0_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product131_1_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product131_1_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product131_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product131_1_impl_out,
                 X => Delay1No170_out_to_Product131_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product131_1_impl_parent_implementedSystem_port_1_cast);

SharedReg175_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg175_out;
Delay3No10_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_2_cast <= Delay3No10_out;
SharedReg189_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg189_out;
SharedReg389_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product131_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg175_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No10_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg189_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product131_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product131_1_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product131_1_impl_0_out,
                 Y => Delay1No170_out);

SharedReg111_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg7_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg391_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product131_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product131_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product131_1_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product131_1_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product131_2_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product131_2_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product131_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product131_2_impl_out,
                 X => Delay1No172_out_to_Product131_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product131_2_impl_parent_implementedSystem_port_1_cast);

SharedReg191_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg389_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg61_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg61_out;
SharedReg61_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg61_out;
   MUX_Product131_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg61_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg61_out_to_MUX_Product131_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product131_2_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product131_2_impl_0_out,
                 Y => Delay1No172_out);

SharedReg391_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg6_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg7_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg7_out;
   MUX_Product131_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg6_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg7_out_to_MUX_Product131_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product131_2_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product131_2_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product371_2_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product371_2_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product371_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product371_2_impl_out,
                 X => Delay1No174_out_to_Product371_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product371_2_impl_parent_implementedSystem_port_1_cast);

SharedReg177_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg177_out;
SharedReg389_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg185_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg185_out;
SharedReg186_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg186_out;
   MUX_Product371_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg177_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg185_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg186_out_to_MUX_Product371_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product371_2_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product371_2_impl_0_out,
                 Y => Delay1No174_out);

SharedReg391_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg21_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg349_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product371_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg21_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product371_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product371_2_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product371_2_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product381_0_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product381_0_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product381_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product381_0_impl_out,
                 X => Delay1No176_out_to_Product381_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product381_0_impl_parent_implementedSystem_port_1_cast);

SharedReg173_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg173_out;
SharedReg172_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg172_out;
SharedReg389_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg180_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg180_out;
   MUX_Product381_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg173_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg172_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg180_out_to_MUX_Product381_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product381_0_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product381_0_impl_0_out,
                 Y => Delay1No176_out);

SharedReg344_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg391_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg114_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
   MUX_Product381_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product381_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product381_0_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product381_0_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product381_1_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product381_1_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product381_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product381_1_impl_out,
                 X => Delay1No178_out_to_Product381_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product381_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
Delay7No58_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_2_cast <= Delay7No58_out;
SharedReg174_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
SharedReg389_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product381_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay7No58_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg174_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product381_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product381_1_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product381_1_impl_0_out,
                 Y => Delay1No178_out);

SharedReg390_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg161_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg391_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product381_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product381_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product381_1_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product381_1_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product391_2_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product391_2_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product391_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product391_2_impl_out,
                 X => Delay1No180_out_to_Product391_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product391_2_impl_parent_implementedSystem_port_1_cast);

SharedReg185_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg185_out;
SharedReg389_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg199_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg199_out;
SharedReg209_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg209_out;
   MUX_Product391_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg185_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg199_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Product391_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product391_2_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product391_2_impl_0_out,
                 Y => Delay1No180_out);

SharedReg391_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg386_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
SharedReg18_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg18_out;
   MUX_Product391_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg18_out_to_MUX_Product391_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product391_2_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product391_2_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product411_0_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product411_0_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product411_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product411_0_impl_out,
                 X => Delay1No182_out_to_Product411_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product411_0_impl_parent_implementedSystem_port_1_cast);

Delay3No15_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No15_out;
SharedReg179_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg179_out;
SharedReg389_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product411_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No15_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg179_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product411_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product411_0_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product411_0_impl_0_out,
                 Y => Delay1No182_out);

SharedReg18_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg391_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product411_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product411_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product411_0_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product411_0_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product411_2_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product411_2_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product411_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product411_2_impl_out,
                 X => Delay1No184_out_to_Product411_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product411_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg214_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg214_out;
   MUX_Product411_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg214_out_to_MUX_Product411_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product411_2_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product411_2_impl_0_out,
                 Y => Delay1No184_out);

SharedReg9_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg12_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg12_out;
   MUX_Product411_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg12_out_to_MUX_Product411_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product411_2_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product411_2_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product421_0_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product421_0_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product421_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product421_0_impl_out,
                 X => Delay1No186_out_to_Product421_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product421_0_impl_parent_implementedSystem_port_1_cast);

SharedReg211_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg211_out;
SharedReg1_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product421_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg211_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product421_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product421_0_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product421_0_impl_0_out,
                 Y => Delay1No186_out);

SharedReg12_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg9_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product421_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product421_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product421_0_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product421_0_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product421_1_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product421_1_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product421_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product421_1_impl_out,
                 X => Delay1No188_out_to_Product421_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product421_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
Delay3No16_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_2_cast <= Delay3No16_out;
SharedReg1_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product421_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No16_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product421_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product421_1_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product421_1_impl_0_out,
                 Y => Delay1No188_out);

SharedReg390_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg18_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg9_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg389_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product421_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product421_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product421_1_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product421_1_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Product421_2_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Product421_2_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Product421_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product421_2_impl_out,
                 X => Delay1No190_out_to_Product421_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Product421_2_impl_parent_implementedSystem_port_1_cast);

SharedReg271_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg271_out;
SharedReg389_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg246_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg246_out;
   MUX_Product421_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg271_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg246_out_to_MUX_Product421_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product421_2_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product421_2_impl_0_out,
                 Y => Delay1No190_out);

SharedReg392_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg389_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg397_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product421_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product421_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product421_2_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product421_2_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Product441_0_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Product441_0_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Product441_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product441_0_impl_out,
                 X => Delay1No192_out_to_Product441_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Product441_0_impl_parent_implementedSystem_port_1_cast);

SharedReg247_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg247_out;
SharedReg274_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg274_out;
SharedReg264_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg264_out;
SharedReg194_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg194_out;
   MUX_Product441_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg247_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg274_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg264_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg194_out_to_MUX_Product441_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product441_0_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_0_impl_0_out,
                 Y => Delay1No192_out);

SharedReg397_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg392_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg396_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg343_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg343_out;
   MUX_Product441_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Product441_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product441_0_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_0_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product441_1_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product441_1_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product441_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product441_1_impl_out,
                 X => Delay1No194_out_to_Product441_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product441_1_impl_parent_implementedSystem_port_1_cast);

SharedReg182_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg206_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg206_out;
SharedReg275_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg275_out;
SharedReg265_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg265_out;
   MUX_Product441_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg206_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg275_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg265_out_to_MUX_Product441_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product441_1_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_1_impl_0_out,
                 Y => Delay1No194_out);

SharedReg160_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg12_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg392_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg396_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product441_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product441_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product441_1_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_1_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Product441_2_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Product441_2_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Product441_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product441_2_impl_out,
                 X => Delay1No196_out_to_Product441_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Product441_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg266_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg266_out;
SharedReg202_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg202_out;
SharedReg219_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg219_out;
   MUX_Product441_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg266_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg202_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg219_out_to_MUX_Product441_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product441_2_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_2_impl_0_out,
                 Y => Delay1No196_out);

SharedReg20_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg396_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg348_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg348_out;
SharedReg22_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg22_out;
   MUX_Product441_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg348_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg22_out_to_MUX_Product441_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product441_2_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product441_2_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product461_0_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product461_0_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product461_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product461_0_impl_out,
                 X => Delay1No198_out_to_Product461_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product461_0_impl_parent_implementedSystem_port_1_cast);

Delay3No21_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No21_out;
SharedReg1_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg215_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg215_out;
   MUX_Product461_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No21_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg215_out_to_MUX_Product461_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product461_0_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_0_impl_0_out,
                 Y => Delay1No198_out);

SharedReg22_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg22_out;
SharedReg20_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg6_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg6_out;
   MUX_Product461_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg22_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg6_out_to_MUX_Product461_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product461_0_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_0_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Product461_1_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Product461_1_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Product461_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product461_1_impl_out,
                 X => Delay1No200_out_to_Product461_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Product461_1_impl_parent_implementedSystem_port_1_cast);

SharedReg216_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg216_out;
SharedReg257_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg257_out;
SharedReg1_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product461_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg216_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product461_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product461_1_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_1_impl_0_out,
                 Y => Delay1No200_out);

SharedReg6_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg6_out;
SharedReg397_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg20_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product461_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product461_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product461_1_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_1_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Product461_2_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Product461_2_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Product461_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product461_2_impl_out,
                 X => Delay1No202_out_to_Product461_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Product461_2_impl_parent_implementedSystem_port_1_cast);

SharedReg227_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg389_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg218_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg218_out;
SharedReg178_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
   MUX_Product461_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg218_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Product461_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product461_2_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_2_impl_0_out,
                 Y => Delay1No202_out);

SharedReg391_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg6_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg12_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg12_out;
   MUX_Product461_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg6_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg12_out_to_MUX_Product461_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product461_2_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product461_2_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Product481_0_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Product481_0_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Product481_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product481_0_impl_out,
                 X => Delay1No204_out_to_Product481_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Product481_0_impl_parent_implementedSystem_port_1_cast);

Delay3No24_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_1_cast <= Delay3No24_out;
SharedReg229_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg229_out;
SharedReg389_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product481_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No24_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product481_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product481_0_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_0_impl_0_out,
                 Y => Delay1No204_out);

SharedReg12_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg12_out;
SharedReg391_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product481_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg12_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product481_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product481_0_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_0_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product481_1_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product481_1_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product481_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product481_1_impl_out,
                 X => Delay1No206_out_to_Product481_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product481_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg217_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg217_out;
SharedReg231_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg231_out;
SharedReg389_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product481_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg217_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg231_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product481_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product481_1_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_1_impl_0_out,
                 Y => Delay1No206_out);

SharedReg390_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg22_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg391_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product481_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product481_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product481_1_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_1_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product481_2_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product481_2_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product481_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product481_2_impl_out,
                 X => Delay1No208_out_to_Product481_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product481_2_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg242_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg242_out;
   MUX_Product481_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg242_out_to_MUX_Product481_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product481_2_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_2_impl_0_out,
                 Y => Delay1No208_out);

SharedReg20_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg390_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg349_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product481_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product481_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product481_2_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product481_2_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product511_0_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product511_0_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product511_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product511_0_impl_out,
                 X => Delay1No210_out_to_Product511_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product511_0_impl_parent_implementedSystem_port_1_cast);

Delay7No60_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_1_cast <= Delay7No60_out;
SharedReg5_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg212_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg212_out;
   MUX_Product511_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay7No60_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg212_out_to_MUX_Product511_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product511_0_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product511_0_impl_0_out,
                 Y => Delay1No210_out);

SharedReg344_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg20_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg105_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product511_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product511_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product511_0_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product511_0_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product511_1_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product511_1_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product511_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product511_1_impl_out,
                 X => Delay1No212_out_to_Product511_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product511_1_impl_parent_implementedSystem_port_1_cast);

Delay5No13_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_1_cast <= Delay5No13_out;
Delay3No25_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_2_cast <= Delay3No25_out;
SharedReg5_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg389_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product511_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No13_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No25_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product511_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product511_1_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product511_1_impl_0_out,
                 Y => Delay1No212_out);

SharedReg169_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg12_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg20_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg389_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product511_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product511_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product511_1_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product511_1_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product511_2_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product511_2_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product511_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product511_2_impl_out,
                 X => Delay1No214_out_to_Product511_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product511_2_impl_parent_implementedSystem_port_1_cast);

SharedReg240_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg240_out;
SharedReg389_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
Delay5No14_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_3_cast <= Delay5No14_out;
SharedReg14_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg14_out;
   MUX_Product511_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg240_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay5No14_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg14_out_to_MUX_Product511_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product511_2_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product511_2_impl_0_out,
                 Y => Delay1No214_out);

SharedReg391_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg351_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg387_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
   MUX_Product511_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg351_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg387_out_to_MUX_Product511_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product511_2_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product511_2_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Product521_0_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Product521_0_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Product521_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product521_0_impl_out,
                 X => Delay1No216_out_to_Product521_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Product521_0_impl_parent_implementedSystem_port_1_cast);

SharedReg14_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg14_out;
SharedReg243_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg243_out;
SharedReg389_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg236_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg236_out;
   MUX_Product521_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg14_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg243_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Product521_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product521_0_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product521_0_impl_0_out,
                 Y => Delay1No216_out);

SharedReg115_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg391_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg105_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product521_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product521_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product521_0_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product521_0_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Product521_1_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Product521_1_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Product521_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product521_1_impl_out,
                 X => Delay1No218_out_to_Product521_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Product521_1_impl_parent_implementedSystem_port_1_cast);

SharedReg238_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg238_out;
SharedReg239_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg239_out;
SharedReg245_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg245_out;
SharedReg389_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product521_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg238_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg239_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg245_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product521_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product521_1_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product521_1_impl_0_out,
                 Y => Delay1No218_out);

SharedReg169_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg161_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg391_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product521_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product521_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product521_1_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product521_1_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Product521_2_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Product521_2_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Product521_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product521_2_impl_out,
                 X => Delay1No220_out_to_Product521_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Product521_2_impl_parent_implementedSystem_port_1_cast);

SharedReg246_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg246_out;
SharedReg389_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg241_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg241_out;
SharedReg322_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg322_out;
   MUX_Product521_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg246_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg241_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg322_out_to_MUX_Product521_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product521_2_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product521_2_impl_0_out,
                 Y => Delay1No220_out);

SharedReg392_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg389_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg351_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg397_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product521_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg351_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product521_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product521_2_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product521_2_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product55_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_0_impl_out,
                 X => Delay1No222_out_to_Product55_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product55_0_impl_parent_implementedSystem_port_1_cast);

Delay2No45_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast <= Delay2No45_out;
SharedReg247_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg247_out;
SharedReg389_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg230_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg230_out;
   MUX_Product55_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No45_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg247_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg230_out_to_MUX_Product55_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_0_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_0_impl_0_out,
                 Y => Delay1No222_out);

SharedReg397_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg392_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg389_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg25_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
   MUX_Product55_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Product55_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_0_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_0_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product55_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_1_impl_out,
                 X => Delay1No224_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast);

SharedReg232_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg232_out;
SharedReg14_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
SharedReg249_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg249_out;
SharedReg389_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product55_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg232_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg249_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_1_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_1_impl_0_out,
                 Y => Delay1No224_out);

SharedReg25_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg112_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg392_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg389_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product55_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_1_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_1_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Product55_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_2_impl_out,
                 X => Delay1No226_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast);

SharedReg24_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg389_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg234_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg234_out;
SharedReg349_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product55_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg234_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_2_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_2_impl_0_out,
                 Y => Delay1No226_out);

SharedReg16_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg25_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg26_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
   MUX_Product55_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_2_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_2_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Product57_0_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Product57_0_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Product57_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product57_0_impl_out,
                 X => Delay1No228_out_to_Product57_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Product57_0_impl_parent_implementedSystem_port_1_cast);

SharedReg344_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg24_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg255_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg255_out;
SharedReg390_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product57_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg255_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product57_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product57_0_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_0_impl_0_out,
                 Y => Delay1No228_out);

SharedReg26_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg16_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg10_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg10_out;
SharedReg390_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product57_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg10_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product57_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product57_0_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_0_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Product57_1_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Product57_1_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Product57_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product57_1_impl_out,
                 X => Delay1No230_out_to_Product57_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Product57_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg320_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg320_out;
SharedReg24_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg257_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg257_out;
   MUX_Product57_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg320_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg257_out_to_MUX_Product57_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product57_1_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_1_impl_0_out,
                 Y => Delay1No230_out);

SharedReg390_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg397_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg16_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg10_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg10_out;
   MUX_Product57_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg10_out_to_MUX_Product57_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product57_1_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_1_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product57_2_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product57_2_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product57_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product57_2_impl_out,
                 X => Delay1No232_out_to_Product57_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product57_2_impl_parent_implementedSystem_port_1_cast);

SharedReg259_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg259_out;
SharedReg259_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg259_out;
SharedReg390_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg4_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg4_out;
   MUX_Product57_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg259_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg259_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg4_out_to_MUX_Product57_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product57_2_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_2_impl_0_out,
                 Y => Delay1No232_out);

SharedReg391_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg10_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg10_out;
SharedReg390_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg387_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
   MUX_Product57_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg10_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg387_out_to_MUX_Product57_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product57_2_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product57_2_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product59_0_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product59_0_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product59_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product59_0_impl_out,
                 X => Delay1No234_out_to_Product59_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product59_0_impl_parent_implementedSystem_port_1_cast);

SharedReg4_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg4_out;
SharedReg260_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg260_out;
SharedReg104_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg390_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product59_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg4_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg260_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product59_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product59_0_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_0_impl_0_out,
                 Y => Delay1No234_out);

SharedReg115_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg391_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg23_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg390_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product59_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg23_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product59_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product59_0_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_0_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Product59_1_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Product59_1_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Product59_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product59_1_impl_out,
                 X => Delay1No236_out_to_Product59_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Product59_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg161_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg261_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg261_out;
SharedReg168_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg168_out;
   MUX_Product59_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg261_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product59_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product59_1_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_1_impl_0_out,
                 Y => Delay1No236_out);

SharedReg390_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg26_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg391_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg23_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg23_out;
   MUX_Product59_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg23_out_to_MUX_Product59_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product59_1_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_1_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Product59_2_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Product59_2_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Product59_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product59_2_impl_out,
                 X => Delay1No238_out_to_Product59_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Product59_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg350_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg390_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg349_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product59_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product59_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product59_2_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_2_impl_0_out,
                 Y => Delay1No238_out);

SharedReg16_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg23_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg390_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg387_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg387_out;
   MUX_Product59_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg387_out_to_MUX_Product59_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product59_2_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product59_2_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Product61_0_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Product61_0_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Product61_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product61_0_impl_out,
                 X => Delay1No240_out_to_Product61_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Product61_0_impl_parent_implementedSystem_port_1_cast);

SharedReg344_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg1_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg260_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg260_out;
   MUX_Product61_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg260_out_to_MUX_Product61_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product61_0_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_0_impl_0_out,
                 Y => Delay1No240_out);

SharedReg115_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg16_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg25_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg25_out;
   MUX_Product61_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg389_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg25_out_to_MUX_Product61_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product61_0_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_0_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Product61_1_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Product61_1_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Product61_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product61_1_impl_out,
                 X => Delay1No242_out_to_Product61_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Product61_1_impl_parent_implementedSystem_port_1_cast);

SharedReg261_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg4_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg1_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg389_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product61_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product61_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product61_1_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_1_impl_0_out,
                 Y => Delay1No242_out);

SharedReg25_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg112_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg16_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg389_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg389_out;
   MUX_Product61_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg389_out_to_MUX_Product61_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product61_1_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_1_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Product61_2_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Product61_2_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Product61_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product61_2_impl_out,
                 X => Delay1No244_out_to_Product61_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Product61_2_impl_parent_implementedSystem_port_1_cast);

SharedReg266_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg389_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg262_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg262_out;
SharedReg259_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg259_out;
   MUX_Product61_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg262_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg259_out_to_MUX_Product61_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product61_2_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_2_impl_0_out,
                 Y => Delay1No244_out);

SharedReg391_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg389_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg389_out;
SharedReg25_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg397_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product61_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg389_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg25_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product61_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product61_2_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product61_2_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product62_0_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product62_0_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product62_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product62_0_impl_out,
                 X => Delay1No246_out_to_Product62_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product62_0_impl_parent_implementedSystem_port_1_cast);

SharedReg260_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg260_out;
SharedReg267_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg267_out;
SharedReg8_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg244_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg244_out;
   MUX_Product62_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg260_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg267_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg8_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_Product62_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product62_0_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_0_impl_0_out,
                 Y => Delay1No246_out);

SharedReg397_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg391_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg104_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg2_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg2_out;
   MUX_Product62_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Product62_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product62_0_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_0_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Product62_1_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Product62_1_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Product62_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product62_1_impl_out,
                 X => Delay1No248_out_to_Product62_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Product62_1_impl_parent_implementedSystem_port_1_cast);

Delay2No43_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_1_cast <= Delay2No43_out;
SharedReg161_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg269_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg269_out;
SharedReg8_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg8_out;
   MUX_Product62_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No43_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg269_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg8_out_to_MUX_Product62_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product62_1_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_1_impl_0_out,
                 Y => Delay1No248_out);

SharedReg2_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg2_out;
SharedReg112_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg391_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg168_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
   MUX_Product62_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product62_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product62_1_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_1_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Product62_2_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Product62_2_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Product62_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product62_2_impl_out,
                 X => Delay1No250_out_to_Product62_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Product62_2_impl_parent_implementedSystem_port_1_cast);

SharedReg233_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg8_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
Delay2No44_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_3_cast <= Delay2No44_out;
SharedReg262_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg262_out;
   MUX_Product62_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No44_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg262_out_to_MUX_Product62_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product62_2_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_2_impl_0_out,
                 Y => Delay1No250_out);

SharedReg392_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg350_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg2_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg397_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product62_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product62_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product62_2_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_2_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Product63_0_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Product63_0_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Product63_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product63_0_impl_out,
                 X => Delay1No252_out_to_Product63_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Product63_0_impl_parent_implementedSystem_port_1_cast);

SharedReg264_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg264_out;
SharedReg235_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg235_out;
SharedReg342_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg342_out;
SharedReg264_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg264_out;
   MUX_Product63_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg264_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg235_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg342_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg264_out_to_MUX_Product63_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product63_0_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_0_impl_0_out,
                 Y => Delay1No252_out);

SharedReg397_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg392_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg104_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg21_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg21_out;
   MUX_Product63_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg21_out_to_MUX_Product63_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product63_0_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_0_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Product63_1_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Product63_1_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Product63_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product63_1_impl_out,
                 X => Delay1No254_out_to_Product63_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Product63_1_impl_parent_implementedSystem_port_1_cast);

SharedReg265_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg265_out;
SharedReg265_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg265_out;
SharedReg237_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg237_out;
SharedReg159_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg159_out;
   MUX_Product63_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg265_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg265_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg237_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product63_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product63_1_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_1_impl_0_out,
                 Y => Delay1No254_out);

SharedReg21_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg21_out;
SharedReg397_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg392_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg168_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
   MUX_Product63_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg21_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product63_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product63_1_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_1_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Product63_2_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Product63_2_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Product63_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product63_2_impl_out,
                 X => Delay1No256_out_to_Product63_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Product63_2_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg347_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg347_out;
SharedReg266_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg266_out;
SharedReg266_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg266_out;
   MUX_Product63_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg347_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg266_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg266_out_to_MUX_Product63_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product63_2_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_2_impl_0_out,
                 Y => Delay1No256_out);

SharedReg9_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg350_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg21_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg21_out;
SharedReg397_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product63_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg21_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product63_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product63_2_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product63_2_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product64_0_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product64_0_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product64_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product64_0_impl_out,
                 X => Delay1No258_out_to_Product64_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product64_0_impl_parent_implementedSystem_port_1_cast);

SharedReg267_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg267_out;
SharedReg5_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg381_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg381_out;
SharedReg390_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product64_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg267_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg381_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product64_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product64_0_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_0_impl_0_out,
                 Y => Delay1No258_out);

SharedReg397_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg9_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg396_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg390_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product64_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product64_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product64_0_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_0_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product64_1_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product64_1_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product64_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product64_1_impl_out,
                 X => Delay1No260_out_to_Product64_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product64_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg269_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg269_out;
SharedReg5_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg382_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg382_out;
   MUX_Product64_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg269_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg382_out_to_MUX_Product64_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product64_1_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_1_impl_0_out,
                 Y => Delay1No260_out);

SharedReg390_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg397_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg9_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg396_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product64_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product64_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product64_1_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_1_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Product64_2_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Product64_2_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Product64_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product64_2_impl_out,
                 X => Delay1No262_out_to_Product64_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Product64_2_impl_parent_implementedSystem_port_1_cast);

SharedReg282_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg282_out;
SharedReg384_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg384_out;
SharedReg390_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg349_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product64_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg282_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg384_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product64_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product64_2_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_2_impl_0_out,
                 Y => Delay1No262_out);

SharedReg391_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg390_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg19_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg19_out;
   MUX_Product64_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg19_out_to_MUX_Product64_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product64_2_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product64_2_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Product66_0_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Product66_0_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Product66_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product66_0_impl_out,
                 X => Delay1No264_out_to_Product66_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Product66_0_impl_parent_implementedSystem_port_1_cast);

SharedReg344_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg283_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg283_out;
SharedReg8_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg390_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product66_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg283_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg8_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product66_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product66_0_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_0_impl_0_out,
                 Y => Delay1No264_out);

SharedReg19_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg391_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg104_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg390_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product66_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product66_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product66_0_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_0_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Product66_1_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Product66_1_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Product66_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product66_1_impl_out,
                 X => Delay1No266_out_to_Product66_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Product66_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg275_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg284_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg284_out;
SharedReg8_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg8_out;
   MUX_Product66_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg284_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg8_out_to_MUX_Product66_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product66_1_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_1_impl_0_out,
                 Y => Delay1No266_out);

SharedReg390_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg397_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg391_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg168_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
   MUX_Product66_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product66_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product66_1_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_1_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Product66_2_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Product66_2_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Product66_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product66_2_impl_out,
                 X => Delay1No268_out_to_Product66_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Product66_2_impl_parent_implementedSystem_port_1_cast);

SharedReg286_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg286_out;
SharedReg8_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg390_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg349_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product66_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg286_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product66_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product66_2_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_2_impl_0_out,
                 Y => Delay1No268_out);

SharedReg392_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg350_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg390_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg19_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg19_out;
   MUX_Product66_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg19_out_to_MUX_Product66_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product66_2_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product66_2_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Product67_0_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Product67_0_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Product67_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product67_0_impl_out,
                 X => Delay1No270_out_to_Product67_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Product67_0_impl_parent_implementedSystem_port_1_cast);

SharedReg344_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg287_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg287_out;
SharedReg287_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg287_out;
SharedReg390_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product67_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg287_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg287_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product67_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product67_0_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_0_impl_0_out,
                 Y => Delay1No270_out);

SharedReg19_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg19_out;
SharedReg392_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg396_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg390_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg390_out;
   MUX_Product67_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg19_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Product67_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product67_0_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_0_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Product67_1_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Product67_1_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Product67_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product67_1_impl_out,
                 X => Delay1No272_out_to_Product67_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Product67_1_impl_parent_implementedSystem_port_1_cast);

SharedReg390_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg161_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg288_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg288_out;
SharedReg288_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg288_out;
   MUX_Product67_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg288_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg288_out_to_MUX_Product67_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product67_1_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_1_impl_0_out,
                 Y => Delay1No272_out);

SharedReg390_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg390_out;
SharedReg19_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg392_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg396_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product67_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg390_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product67_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product67_1_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_1_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Product67_2_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Product67_2_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Product67_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product67_2_impl_out,
                 X => Delay1No274_out_to_Product67_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Product67_2_impl_parent_implementedSystem_port_1_cast);

SharedReg5_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg5_out;
SharedReg289_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg289_out;
SharedReg390_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg289_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg289_out;
   MUX_Product67_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg5_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg289_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg289_out_to_MUX_Product67_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product67_2_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_2_impl_0_out,
                 Y => Delay1No274_out);

SharedReg24_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg396_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg390_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg390_out;
SharedReg397_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product67_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg390_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product67_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product67_2_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_2_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Product68_0_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Product68_0_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Product68_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product68_0_impl_out,
                 X => Delay1No276_out_to_Product68_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Product68_0_impl_parent_implementedSystem_port_1_cast);

SharedReg291_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg291_out;
SharedReg5_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg113_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg113_out;
SharedReg283_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg283_out;
   MUX_Product68_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg113_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg283_out_to_MUX_Product68_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product68_0_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_0_impl_0_out,
                 Y => Delay1No276_out);

SharedReg397_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg24_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg13_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg13_out;
SharedReg2_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg2_out;
   MUX_Product68_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg13_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Product68_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product68_0_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_0_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Product68_1_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Product68_1_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Product68_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product68_1_impl_out,
                 X => Delay1No278_out_to_Product68_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Product68_1_impl_parent_implementedSystem_port_1_cast);

SharedReg284_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg284_out;
SharedReg161_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg5_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg5_out;
SharedReg110_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg110_out;
   MUX_Product68_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg284_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg5_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Product68_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product68_1_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_1_impl_0_out,
                 Y => Delay1No278_out);

SharedReg2_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg2_out;
SharedReg19_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg24_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg13_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg13_out;
   MUX_Product68_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg13_out_to_MUX_Product68_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product68_1_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_1_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Product68_2_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Product68_2_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Product68_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product68_2_impl_out,
                 X => Delay1No280_out_to_Product68_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Product68_2_impl_parent_implementedSystem_port_1_cast);

SharedReg297_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg297_out;
SharedReg385_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg385_out;
SharedReg286_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg286_out;
SharedReg297_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg297_out;
   MUX_Product68_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg297_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg385_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg286_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg297_out_to_MUX_Product68_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product68_2_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_2_impl_0_out,
                 Y => Delay1No280_out);

SharedReg391_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg13_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg2_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg400_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
   MUX_Product68_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Product68_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product68_2_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_2_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Product711_0_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Product711_0_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Product711_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product711_0_impl_out,
                 X => Delay1No282_out_to_Product711_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Product711_0_impl_parent_implementedSystem_port_1_cast);

SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg299_out;
SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg299_out;
SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg299_out;
SharedReg248_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg248_out;
   MUX_Product711_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg299_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg248_out_to_MUX_Product711_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product711_0_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product711_0_impl_0_out,
                 Y => Delay1No282_out);

SharedReg400_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg400_out;
SharedReg391_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg114_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
   MUX_Product711_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product711_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product711_0_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product711_0_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Product711_1_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Product711_1_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Product711_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product711_1_impl_out,
                 X => Delay1No284_out_to_Product711_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Product711_1_impl_parent_implementedSystem_port_1_cast);

SharedReg250_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg250_out;
SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg300_out;
SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg300_out;
   MUX_Product711_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg250_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg300_out_to_MUX_Product711_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product711_1_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product711_1_impl_0_out,
                 Y => Delay1No284_out);

SharedReg111_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg397_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg391_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product711_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product711_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product711_1_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product711_1_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Product711_2_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Product711_2_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Product711_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product711_2_impl_out,
                 X => Delay1No286_out_to_Product711_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Product711_2_impl_parent_implementedSystem_port_1_cast);

SharedReg24_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg24_out;
SharedReg301_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg301_out;
SharedReg253_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg253_out;
SharedReg380_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg380_out;
   MUX_Product711_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg24_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg301_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg253_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg380_out_to_MUX_Product711_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product711_2_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product711_2_impl_0_out,
                 Y => Delay1No286_out);

SharedReg9_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg396_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg386_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
SharedReg397_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product711_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product711_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product711_2_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product711_2_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Product70_0_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Product70_0_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Product70_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product70_0_impl_out,
                 X => Delay1No288_out_to_Product70_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Product70_0_impl_parent_implementedSystem_port_1_cast);

SharedReg375_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg375_out;
SharedReg24_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg304_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg304_out;
Delay5No18_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_4_cast <= Delay5No18_out;
   MUX_Product70_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg375_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg304_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No18_out_to_MUX_Product70_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product70_0_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_0_impl_0_out,
                 Y => Delay1No288_out);

SharedReg397_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg9_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg398_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg398_out;
SharedReg343_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg343_out;
   MUX_Product70_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg398_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Product70_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product70_0_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_0_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Product70_1_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Product70_1_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Product70_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product70_1_impl_out,
                 X => Delay1No290_out_to_Product70_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Product70_1_impl_parent_implementedSystem_port_1_cast);

Delay5No19_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_1_cast <= Delay5No19_out;
SharedReg306_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg306_out;
SharedReg24_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg306_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg306_out;
   MUX_Product70_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No19_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg306_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg24_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg306_out_to_MUX_Product70_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product70_1_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_1_impl_0_out,
                 Y => Delay1No290_out);

SharedReg160_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg400_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg400_out;
SharedReg9_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg398_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg398_out;
   MUX_Product70_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg400_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg398_out_to_MUX_Product70_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product70_1_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_1_impl_1_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Product70_2_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Product70_2_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Product70_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product70_2_impl_out,
                 X => Delay1No292_out_to_Product70_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Product70_2_impl_parent_implementedSystem_port_1_cast);

SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg307_out;
SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg307_out;
SharedReg290_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg290_out;
SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg307_out;
   MUX_Product70_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg290_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg307_out_to_MUX_Product70_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product70_2_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_2_impl_0_out,
                 Y => Delay1No292_out);

SharedReg391_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg398_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg398_out;
SharedReg348_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg348_out;
SharedReg400_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
   MUX_Product70_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg398_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg348_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Product70_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product70_2_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product70_2_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Product71_0_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Product71_0_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Product71_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product71_0_impl_out,
                 X => Delay1No294_out_to_Product71_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Product71_0_impl_parent_implementedSystem_port_1_cast);

SharedReg308_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg308_out;
SharedReg308_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg308_out;
SharedReg23_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg293_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg293_out;
   MUX_Product71_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg308_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg308_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg23_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg293_out_to_MUX_Product71_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product71_0_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_0_impl_0_out,
                 Y => Delay1No294_out);

SharedReg400_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg400_out;
SharedReg391_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg104_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg105_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product71_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product71_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product71_0_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_0_impl_1_out,
                 Y => Delay1No295_out);

Delay1No296_out_to_Product71_1_impl_parent_implementedSystem_port_0_cast <= Delay1No296_out;
Delay1No297_out_to_Product71_1_impl_parent_implementedSystem_port_1_cast <= Delay1No297_out;
   Product71_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product71_1_impl_out,
                 X => Delay1No296_out_to_Product71_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No297_out_to_Product71_1_impl_parent_implementedSystem_port_1_cast);

SharedReg296_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg296_out;
SharedReg378_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg378_out;
SharedReg309_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg309_out;
SharedReg23_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg23_out;
   MUX_Product71_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg296_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg378_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg309_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg23_out_to_MUX_Product71_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product71_1_impl_0_out);

   Delay1No296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_1_impl_0_out,
                 Y => Delay1No296_out);

SharedReg169_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg397_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg391_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg168_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg168_out;
   MUX_Product71_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg168_out_to_MUX_Product71_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product71_1_impl_1_out);

   Delay1No297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_1_impl_1_out,
                 Y => Delay1No297_out);

Delay1No298_out_to_Product71_2_impl_parent_implementedSystem_port_0_cast <= Delay1No298_out;
Delay1No299_out_to_Product71_2_impl_parent_implementedSystem_port_1_cast <= Delay1No299_out;
   Product71_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product71_2_impl_out,
                 X => Delay1No298_out_to_Product71_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No299_out_to_Product71_2_impl_parent_implementedSystem_port_1_cast);

SharedReg20_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg20_out;
SharedReg23_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg23_out;
Delay5No23_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_3_cast <= Delay5No23_out;
SharedReg349_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg349_out;
   MUX_Product71_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg20_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay5No23_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg349_out_to_MUX_Product71_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product71_2_impl_0_out);

   Delay1No298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_2_impl_0_out,
                 Y => Delay1No298_out);

SharedReg16_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg16_out;
SharedReg350_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg351_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg26_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg26_out;
   MUX_Product71_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg16_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg351_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Product71_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product71_2_impl_1_out);

   Delay1No299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product71_2_impl_1_out,
                 Y => Delay1No299_out);

Delay1No300_out_to_Product76_0_impl_parent_implementedSystem_port_0_cast <= Delay1No300_out;
Delay1No301_out_to_Product76_0_impl_parent_implementedSystem_port_1_cast <= Delay1No301_out;
   Product76_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product76_0_impl_out,
                 X => Delay1No300_out_to_Product76_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No301_out_to_Product76_0_impl_parent_implementedSystem_port_1_cast);

SharedReg344_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg344_out;
SharedReg20_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg314_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg314_out;
SharedReg105_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product76_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg344_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg314_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product76_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product76_0_impl_0_out);

   Delay1No300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_0_impl_0_out,
                 Y => Delay1No300_out);

SharedReg26_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg16_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg396_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg114_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg114_out;
   MUX_Product76_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product76_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product76_0_impl_1_out);

   Delay1No301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_0_impl_1_out,
                 Y => Delay1No301_out);

Delay1No302_out_to_Product76_1_impl_parent_implementedSystem_port_0_cast <= Delay1No302_out;
Delay1No303_out_to_Product76_1_impl_parent_implementedSystem_port_1_cast <= Delay1No303_out;
   Product76_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product76_1_impl_out,
                 X => Delay1No302_out_to_Product76_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No303_out_to_Product76_1_impl_parent_implementedSystem_port_1_cast);

SharedReg169_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg316_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg316_out;
SharedReg20_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg20_out;
SharedReg316_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg316_out;
   MUX_Product76_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg316_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg20_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg316_out_to_MUX_Product76_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product76_1_impl_0_out);

   Delay1No302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_1_impl_0_out,
                 Y => Delay1No302_out);

SharedReg111_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg400_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg400_out;
SharedReg16_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg16_out;
SharedReg396_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product76_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg400_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg16_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product76_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product76_1_impl_1_out);

   Delay1No303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_1_impl_1_out,
                 Y => Delay1No303_out);

Delay1No304_out_to_Product76_2_impl_parent_implementedSystem_port_0_cast <= Delay1No304_out;
Delay1No305_out_to_Product76_2_impl_parent_implementedSystem_port_1_cast <= Delay1No305_out;
   Product76_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product76_2_impl_out,
                 X => Delay1No304_out_to_Product76_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No305_out_to_Product76_2_impl_parent_implementedSystem_port_1_cast);

SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg351_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg317_out;
   MUX_Product76_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg351_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg317_out_to_MUX_Product76_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product76_2_impl_0_out);

   Delay1No304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_2_impl_0_out,
                 Y => Delay1No304_out);

SharedReg391_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg386_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
SharedReg397_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product76_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product76_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product76_2_impl_1_out);

   Delay1No305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product76_2_impl_1_out,
                 Y => Delay1No305_out);

Delay1No306_out_to_Product911_0_impl_parent_implementedSystem_port_0_cast <= Delay1No306_out;
Delay1No307_out_to_Product911_0_impl_parent_implementedSystem_port_1_cast <= Delay1No307_out;
   Product911_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product911_0_impl_out,
                 X => Delay1No306_out_to_Product911_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No307_out_to_Product911_0_impl_parent_implementedSystem_port_1_cast);

SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg318_out;
SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg318_out;
SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg318_out;
SharedReg268_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg268_out;
   MUX_Product911_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg318_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg268_out_to_MUX_Product911_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product911_0_impl_0_out);

   Delay1No306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_0_impl_0_out,
                 Y => Delay1No306_out);

SharedReg397_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg391_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg398_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg398_out;
SharedReg2_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg2_out;
   MUX_Product911_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg398_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg2_out_to_MUX_Product911_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product911_0_impl_1_out);

   Delay1No307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_0_impl_1_out,
                 Y => Delay1No307_out);

Delay1No308_out_to_Product911_1_impl_parent_implementedSystem_port_0_cast <= Delay1No308_out;
Delay1No309_out_to_Product911_1_impl_parent_implementedSystem_port_1_cast <= Delay1No309_out;
   Product911_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product911_1_impl_out,
                 X => Delay1No308_out_to_Product911_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No309_out_to_Product911_1_impl_parent_implementedSystem_port_1_cast);

SharedReg270_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg270_out;
SharedReg161_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg161_out;
SharedReg319_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg319_out;
SharedReg319_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg319_out;
   MUX_Product911_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg270_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg161_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg319_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg319_out_to_MUX_Product911_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product911_1_impl_0_out);

   Delay1No308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_1_impl_0_out,
                 Y => Delay1No308_out);

SharedReg2_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg2_out;
SharedReg26_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg26_out;
SharedReg391_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg398_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg398_out;
   MUX_Product911_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg2_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg26_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg398_out_to_MUX_Product911_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product911_1_impl_1_out);

   Delay1No309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_1_impl_1_out,
                 Y => Delay1No309_out);

Delay1No310_out_to_Product911_2_impl_parent_implementedSystem_port_0_cast <= Delay1No310_out;
Delay1No311_out_to_Product911_2_impl_parent_implementedSystem_port_1_cast <= Delay1No311_out;
   Product911_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product911_2_impl_out,
                 X => Delay1No310_out_to_Product911_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No311_out_to_Product911_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1_out;
SharedReg321_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg321_out;
SharedReg272_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg272_out;
SharedReg302_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg302_out;
   MUX_Product911_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg321_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg272_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg302_out_to_MUX_Product911_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product911_2_impl_0_out);

   Delay1No310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_2_impl_0_out,
                 Y => Delay1No310_out);

SharedReg9_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg9_out;
SharedReg398_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg398_out;
SharedReg2_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg2_out;
SharedReg395_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg395_out;
   MUX_Product911_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg9_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg398_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg2_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg395_out_to_MUX_Product911_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product911_2_impl_1_out);

   Delay1No311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product911_2_impl_1_out,
                 Y => Delay1No311_out);

Delay1No312_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No312_out;
Delay1No313_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No313_out;
   Subtract12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_0_impl_out,
                 X => Delay1No312_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No313_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg87_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg87_out;
SharedReg188_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg188_out;
Delay18No3_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast <= Delay18No3_out;
SharedReg43_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg43_out;
   MUX_Subtract12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg87_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg188_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay18No3_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg43_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract12_0_impl_0_out);

   Delay1No312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_0_out,
                 Y => Delay1No312_out);

SharedReg99_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg134_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg134_out;
SharedReg147_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg147_out;
SharedReg120_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg120_out;
   MUX_Subtract12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg134_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg147_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg120_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract12_0_impl_1_out);

   Delay1No313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_1_out,
                 Y => Delay1No313_out);

Delay1No314_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No314_out;
Delay1No315_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No315_out;
   Subtract12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_1_impl_out,
                 X => Delay1No314_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No315_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast);

Delay11No9_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast <= Delay11No9_out;
SharedReg81_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg81_out;
SharedReg190_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg190_out;
Delay18No4_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast <= Delay18No4_out;
   MUX_Subtract12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No9_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg190_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay18No4_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract12_1_impl_0_out);

   Delay1No314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_0_out,
                 Y => Delay1No314_out);

SharedReg130_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg130_out;
SharedReg101_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg101_out;
SharedReg135_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg135_out;
Delay2No1_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast <= Delay2No1_out;
   MUX_Subtract12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg130_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg135_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No1_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract12_1_impl_1_out);

   Delay1No315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_1_out,
                 Y => Delay1No315_out);

Delay1No316_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No316_out;
Delay1No317_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No317_out;
   Subtract12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_2_impl_out,
                 X => Delay1No316_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No317_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg370_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg370_out;
Delay11No10_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast <= Delay11No10_out;
Delay6No5_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast <= Delay6No5_out;
SharedReg98_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg98_out;
   MUX_Subtract12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg370_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay11No10_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay6No5_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg98_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract12_2_impl_0_out);

   Delay1No316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_0_out,
                 Y => Delay1No316_out);

Delay4No7_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast <= Delay4No7_out;
SharedReg132_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
SharedReg133_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg133_out;
SharedReg102_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg102_out;
   MUX_Subtract12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay4No7_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg133_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg102_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract12_2_impl_1_out);

   Delay1No317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_1_out,
                 Y => Delay1No317_out);

Delay1No318_out_to_Subtract1_2_impl_parent_implementedSystem_port_0_cast <= Delay1No318_out;
Delay1No319_out_to_Subtract1_2_impl_parent_implementedSystem_port_1_cast <= Delay1No319_out;
   Subtract1_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract1_2_impl_out,
                 X => Delay1No318_out_to_Subtract1_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No319_out_to_Subtract1_2_impl_parent_implementedSystem_port_1_cast);

SharedReg192_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg192_out;
Delay18No5_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_2_cast <= Delay18No5_out;
SharedReg228_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg228_out;
SharedReg65_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg65_out;
   MUX_Subtract1_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg192_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay18No5_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg228_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg65_out_to_MUX_Subtract1_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract1_2_impl_0_out);

   Delay1No318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_2_impl_0_out,
                 Y => Delay1No318_out);

SharedReg133_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg151_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg151_out;
SharedReg103_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg156_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg156_out;
   MUX_Subtract1_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg151_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg156_out_to_MUX_Subtract1_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract1_2_impl_1_out);

   Delay1No319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract1_2_impl_1_out,
                 Y => Delay1No319_out);

Delay1No320_out_to_Subtract11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No320_out;
Delay1No321_out_to_Subtract11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No321_out;
   Subtract11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract11_1_impl_out,
                 X => Delay1No320_out_to_Subtract11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No321_out_to_Subtract11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg38_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg53_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg183_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg183_out;
Delay8No28_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_4_cast <= Delay8No28_out;
   MUX_Subtract11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg183_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay8No28_out_to_MUX_Subtract11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract11_1_impl_0_out);

   Delay1No320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_1_impl_0_out,
                 Y => Delay1No320_out);

SharedReg101_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg149_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg149_out;
SharedReg168_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg122_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg122_out;
   MUX_Subtract11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg168_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_Subtract11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract11_1_impl_1_out);

   Delay1No321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_1_impl_1_out,
                 Y => Delay1No321_out);

Delay1No322_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No322_out;
Delay1No323_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No323_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No322_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No323_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg57_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg57_out;
SharedReg195_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg195_out;
Delay8No27_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= Delay8No27_out;
Delay8No21_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= Delay8No21_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg57_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg195_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay8No27_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay8No21_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No322_out);

SharedReg146_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg146_out;
SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg167_out;
SharedReg121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg121_out;
SharedReg121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg121_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg146_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg167_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg121_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No323_out);

Delay1No324_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No324_out;
Delay1No325_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No325_out;
   Subtract3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_0_impl_out,
                 X => Delay1No324_out_to_Subtract3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No325_out_to_Subtract3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg32_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
Delay6No18_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast <= Delay6No18_out;
Delay22No_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast <= Delay22No_out;
SharedReg367_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg367_out;
   MUX_Subtract3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay6No18_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg367_out_to_MUX_Subtract3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_0_impl_0_out);

   Delay1No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_0_out,
                 Y => Delay1No324_out);

SharedReg153_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg99_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg99_out;
SharedReg124_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg124_out;
SharedReg106_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg106_out;
   MUX_Subtract3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg99_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg124_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg106_out_to_MUX_Subtract3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_0_impl_1_out);

   Delay1No325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_0_impl_1_out,
                 Y => Delay1No325_out);

Delay1No326_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No326_out;
Delay1No327_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No327_out;
   Subtract3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_1_impl_out,
                 X => Delay1No326_out_to_Subtract3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No327_out_to_Subtract3_1_impl_parent_implementedSystem_port_1_cast);

Delay8No22_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast <= Delay8No22_out;
SharedReg171_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg171_out;
Delay6No19_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast <= Delay6No19_out;
Delay22No1_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast <= Delay22No1_out;
   MUX_Subtract3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay8No22_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg171_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay6No19_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay22No1_out_to_MUX_Subtract3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_1_impl_0_out);

   Delay1No326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_0_out,
                 Y => Delay1No326_out);

SharedReg122_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg155_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg155_out;
SharedReg101_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg101_out;
SharedReg101_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg101_out;
   MUX_Subtract3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg155_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg101_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Subtract3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_1_impl_1_out);

   Delay1No327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_1_impl_1_out,
                 Y => Delay1No327_out);

Delay1No328_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No328_out;
Delay1No329_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No329_out;
   Subtract3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_2_impl_out,
                 X => Delay1No328_out_to_Subtract3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No329_out_to_Subtract3_2_impl_parent_implementedSystem_port_1_cast);

Delay11No8_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast <= Delay11No8_out;
SharedReg273_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg273_out;
SharedReg373_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg373_out;
SharedReg40_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg40_out;
   MUX_Subtract3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay11No8_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg273_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg373_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg40_out_to_MUX_Subtract3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_2_impl_0_out);

   Delay1No328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_2_impl_0_out,
                 Y => Delay1No328_out);

SharedReg164_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg108_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg108_out;
Delay4No8_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast <= Delay4No8_out;
SharedReg162_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg162_out;
   MUX_Subtract3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay4No8_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg162_out_to_MUX_Subtract3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_2_impl_1_out);

   Delay1No329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_2_impl_1_out,
                 Y => Delay1No329_out);

Delay1No330_out_to_Subtract5_2_impl_parent_implementedSystem_port_0_cast <= Delay1No330_out;
Delay1No331_out_to_Subtract5_2_impl_parent_implementedSystem_port_1_cast <= Delay1No331_out;
   Subtract5_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract5_2_impl_out,
                 X => Delay1No330_out_to_Subtract5_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No331_out_to_Subtract5_2_impl_parent_implementedSystem_port_1_cast);

Delay6No20_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_1_cast <= Delay6No20_out;
Delay11No11_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_2_cast <= Delay11No11_out;
Delay22No2_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_3_cast <= Delay22No2_out;
   MUX_Subtract5_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay6No20_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay11No11_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No2_out_to_MUX_Subtract5_2_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Subtract5_2_impl_0_LUT_out,
                 oMux => MUX_Subtract5_2_impl_0_out);

   Delay1No330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_2_impl_0_out,
                 Y => Delay1No330_out);

SharedReg110_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg133_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg133_out;
SharedReg133_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg133_out;
   MUX_Subtract5_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg133_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg133_out_to_MUX_Subtract5_2_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Subtract5_2_impl_1_LUT_out,
                 oMux => MUX_Subtract5_2_impl_1_out);

   Delay1No331_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract5_2_impl_1_out,
                 Y => Delay1No331_out);

Delay1No332_out_to_Add32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No332_out;
Delay1No333_out_to_Add32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No333_out;
   Add32_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add32_0_impl_out,
                 X => Delay1No332_out_to_Add32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No333_out_to_Add32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg381_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg381_out;
SharedReg_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
Delay57No_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_3_cast <= Delay57No_out;
Delay27No_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_4_cast <= Delay27No_out;
   MUX_Add32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg381_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay57No_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay27No_out_to_MUX_Add32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add32_0_impl_0_out);

   Delay1No332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add32_0_impl_0_out,
                 Y => Delay1No332_out);

SharedReg376_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg376_out;
SharedReg374_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg374_out;
SharedReg114_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg114_out;
SharedReg158_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg158_out;
   MUX_Add32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg376_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg374_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg114_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg158_out_to_MUX_Add32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add32_0_impl_1_out);

   Delay1No333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add32_0_impl_1_out,
                 Y => Delay1No333_out);

Delay1No334_out_to_Add32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No334_out;
Delay1No335_out_to_Add32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No335_out;
   Add32_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add32_2_impl_out,
                 X => Delay1No334_out_to_Add32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No335_out_to_Add32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg358_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg358_out;
Delay95No2_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_2_cast <= Delay95No2_out;
Delay73No2_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_3_cast <= Delay73No2_out;
SharedReg379_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg379_out;
   MUX_Add32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg358_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay95No2_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay73No2_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Add32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add32_2_impl_0_out);

   Delay1No334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add32_2_impl_0_out,
                 Y => Delay1No334_out);

SharedReg345_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg345_out;
SharedReg166_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg166_out;
SharedReg156_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg156_out;
Delay11No14_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_4_cast <= Delay11No14_out;
   MUX_Add32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg345_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg166_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg156_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay11No14_out_to_MUX_Add32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add32_2_impl_1_out);

   Delay1No335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add32_2_impl_1_out,
                 Y => Delay1No335_out);

Delay1No336_out_to_Add211_2_impl_parent_implementedSystem_port_0_cast <= Delay1No336_out;
Delay1No337_out_to_Add211_2_impl_parent_implementedSystem_port_1_cast <= Delay1No337_out;
   Add211_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add211_2_impl_out,
                 X => Delay1No336_out_to_Add211_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No337_out_to_Add211_2_impl_parent_implementedSystem_port_1_cast);

Delay37No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_1_cast <= Delay37No2_out;
SharedReg331_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg331_out;
Delay27No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_3_cast <= Delay27No2_out;
Delay32No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_4_cast <= Delay32No2_out;
   MUX_Add211_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay37No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg331_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay27No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay32No2_out_to_MUX_Add211_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add211_2_impl_0_out);

   Delay1No336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add211_2_impl_0_out,
                 Y => Delay1No336_out);

SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg345_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg346_out;
SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg346_out;
   MUX_Add211_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg346_out_to_MUX_Add211_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add211_2_impl_1_out);

   Delay1No337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add211_2_impl_1_out,
                 Y => Delay1No337_out);

Delay1No338_out_to_Add6_2_impl_parent_implementedSystem_port_0_cast <= Delay1No338_out;
Delay1No339_out_to_Add6_2_impl_parent_implementedSystem_port_1_cast <= Delay1No339_out;
   Add6_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add6_2_impl_out,
                 X => Delay1No338_out_to_Add6_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No339_out_to_Add6_2_impl_parent_implementedSystem_port_1_cast);

SharedReg_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg_out;
SharedReg372_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg313_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg313_out;
Delay51No2_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_4_cast <= Delay51No2_out;
   MUX_Add6_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg313_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay51No2_out_to_MUX_Add6_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add6_2_impl_0_out);

   Delay1No338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_2_impl_0_out,
                 Y => Delay1No338_out);

SharedReg371_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg371_out;
SharedReg346_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg347_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg347_out;
SharedReg340_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg340_out;
   MUX_Add6_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg371_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg347_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg340_out_to_MUX_Add6_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add6_2_impl_1_out);

   Delay1No339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_2_impl_1_out,
                 Y => Delay1No339_out);

Delay1No340_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No340_out;
Delay1No341_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No341_out;
   Add9_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_2_impl_out,
                 X => Delay1No340_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No341_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg15_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg15_out;
Delay57No2_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast <= Delay57No2_out;
   MUX_Add9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg15_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay57No2_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add9_2_impl_0_LUT_out,
                 oMux => MUX_Add9_2_impl_0_out);

   Delay1No340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_2_impl_0_out,
                 Y => Delay1No340_out);

SharedReg348_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg379_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg379_out;
   MUX_Add9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg379_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add9_2_impl_1_LUT_out,
                 oMux => MUX_Add9_2_impl_1_out);

   Delay1No341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_2_impl_1_out,
                 Y => Delay1No341_out);
   Constant1_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

Delay1No342_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast <= Delay1No342_out;
Delay1No343_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast <= Delay1No343_out;
   Divide_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_0_impl_out,
                 X => Delay1No342_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No343_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast);

SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg352_out;
SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg352_out;
SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg352_out;
   MUX_Divide_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg352_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Divide_0_impl_0_LUT_out,
                 oMux => MUX_Divide_0_impl_0_out);

   Delay1No342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_0_out,
                 Y => Delay1No342_out);

SharedReg153_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg153_out;
SharedReg149_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg149_out;
SharedReg345_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg345_out;
   MUX_Divide_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg153_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg345_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Divide_0_impl_1_LUT_out,
                 oMux => MUX_Divide_0_impl_1_out);

   Delay1No343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_1_out,
                 Y => Delay1No343_out);

Delay1No344_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No344_out;
Delay1No345_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No345_out;
   Product11_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_0_impl_out,
                 X => Delay1No344_out_to_Product11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No345_out_to_Product11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg305_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg305_out;
SharedReg1_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg342_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg342_out;
Delay2No54_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast <= Delay2No54_out;
   MUX_Product11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg305_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg342_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No54_out_to_MUX_Product11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_0_impl_0_out);

   Delay1No344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_0_impl_0_out,
                 Y => Delay1No344_out);

SharedReg395_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg395_out;
SharedReg9_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg113_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg113_out;
SharedReg399_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg399_out;
   MUX_Product11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg395_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg113_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg399_out_to_MUX_Product11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_0_impl_1_out);

   Delay1No345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_0_impl_1_out,
                 Y => Delay1No345_out);

Delay1No346_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No346_out;
Delay1No347_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No347_out;
   Product11_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_1_impl_out,
                 X => Delay1No346_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No347_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg285_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg285_out;
SharedReg326_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg326_out;
SharedReg1_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg159_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg159_out;
   MUX_Product11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg285_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg326_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_1_impl_0_out);

   Delay1No346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_0_out,
                 Y => Delay1No346_out);

SharedReg399_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg399_out;
SharedReg397_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg9_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg110_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg110_out;
   MUX_Product11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg399_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg9_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_1_impl_1_out);

   Delay1No347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_1_out,
                 Y => Delay1No347_out);

Delay1No348_out_to_Product11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No348_out;
Delay1No349_out_to_Product11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No349_out;
   Product11_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_2_impl_out,
                 X => Delay1No348_out_to_Product11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No349_out_to_Product11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg329_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg329_out;
SharedReg347_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg347_out;
Delay2No56_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_3_cast <= Delay2No56_out;
SharedReg312_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg312_out;
   MUX_Product11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg329_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg347_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No56_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg312_out_to_MUX_Product11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_2_impl_0_out);

   Delay1No348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_2_impl_0_out,
                 Y => Delay1No348_out);

SharedReg391_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg385_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg385_out;
SharedReg399_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg399_out;
SharedReg395_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg395_out;
   MUX_Product11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg385_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg399_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg395_out_to_MUX_Product11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_2_impl_1_out);

   Delay1No349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_2_impl_1_out,
                 Y => Delay1No349_out);

Delay1No350_out_to_Product14_0_impl_parent_implementedSystem_port_0_cast <= Delay1No350_out;
Delay1No351_out_to_Product14_0_impl_parent_implementedSystem_port_1_cast <= Delay1No351_out;
   Product14_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product14_0_impl_out,
                 X => Delay1No350_out_to_Product14_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No351_out_to_Product14_0_impl_parent_implementedSystem_port_1_cast);

SharedReg315_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg315_out;
SharedReg354_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg354_out;
SharedReg354_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg354_out;
SharedReg292_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg292_out;
   MUX_Product14_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg315_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg354_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg354_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg292_out_to_MUX_Product14_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product14_0_impl_0_out);

   Delay1No350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_0_impl_0_out,
                 Y => Delay1No350_out);

SharedReg395_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg395_out;
SharedReg391_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg399_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg399_out;
   MUX_Product14_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg395_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg396_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg399_out_to_MUX_Product14_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product14_0_impl_1_out);

   Delay1No351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_0_impl_1_out,
                 Y => Delay1No351_out);

Delay1No352_out_to_Product14_1_impl_parent_implementedSystem_port_0_cast <= Delay1No352_out;
Delay1No353_out_to_Product14_1_impl_parent_implementedSystem_port_1_cast <= Delay1No353_out;
   Product14_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product14_1_impl_out,
                 X => Delay1No352_out_to_Product14_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No353_out_to_Product14_1_impl_parent_implementedSystem_port_1_cast);

SharedReg295_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg295_out;
Delay4No46_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No46_out;
SharedReg356_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg356_out;
SharedReg356_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg356_out;
   MUX_Product14_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg295_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No46_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg356_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg356_out_to_MUX_Product14_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product14_1_impl_0_out);

   Delay1No352_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_1_impl_0_out,
                 Y => Delay1No352_out);

SharedReg399_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg399_out;
SharedReg395_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg395_out;
SharedReg391_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg391_out;
SharedReg396_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg396_out;
   MUX_Product14_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg399_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg395_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg391_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg396_out_to_MUX_Product14_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product14_1_impl_1_out);

   Delay1No353_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_1_impl_1_out,
                 Y => Delay1No353_out);

Delay1No354_out_to_Product14_2_impl_parent_implementedSystem_port_0_cast <= Delay1No354_out;
Delay1No355_out_to_Product14_2_impl_parent_implementedSystem_port_1_cast <= Delay1No355_out;
   Product14_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product14_2_impl_out,
                 X => Delay1No354_out_to_Product14_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No355_out_to_Product14_2_impl_parent_implementedSystem_port_1_cast);

SharedReg357_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg357_out;
SharedReg357_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg357_out;
SharedReg298_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg298_out;
Delay2No65_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_4_cast <= Delay2No65_out;
   MUX_Product14_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg357_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg357_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg298_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No65_out_to_MUX_Product14_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product14_2_impl_0_out);

   Delay1No354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_2_impl_0_out,
                 Y => Delay1No354_out);

SharedReg392_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg396_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg399_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg399_out;
SharedReg397_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg397_out;
   MUX_Product14_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg399_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Product14_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product14_2_impl_1_out);

   Delay1No355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product14_2_impl_1_out,
                 Y => Delay1No355_out);

Delay1No356_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast <= Delay1No356_out;
Delay1No357_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast <= Delay1No357_out;
   Product26_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_0_impl_out,
                 X => Delay1No356_out_to_Product26_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No357_out_to_Product26_0_impl_parent_implementedSystem_port_1_cast);

Delay2No63_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast <= Delay2No63_out;
SharedReg359_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg359_out;
SharedReg359_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg359_out;
Delay3No33_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast <= Delay3No33_out;
   MUX_Product26_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No63_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg359_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg359_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No33_out_to_MUX_Product26_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product26_0_impl_0_out);

   Delay1No356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_0_out,
                 Y => Delay1No356_out);

SharedReg397_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg397_out;
SharedReg392_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg392_out;
SharedReg398_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg398_out;
SharedReg394_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg394_out;
   MUX_Product26_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg397_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg392_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg398_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg394_out_to_MUX_Product26_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product26_0_impl_1_out);

   Delay1No357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_0_impl_1_out,
                 Y => Delay1No357_out);

Delay1No358_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No358_out;
Delay1No359_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No359_out;
   Product26_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_1_impl_out,
                 X => Delay1No358_out_to_Product26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No359_out_to_Product26_1_impl_parent_implementedSystem_port_1_cast);

Delay3No34_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast <= Delay3No34_out;
Delay4No49_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast <= Delay4No49_out;
SharedReg361_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg361_out;
SharedReg361_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg361_out;
   MUX_Product26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No34_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No49_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg361_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg361_out_to_MUX_Product26_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product26_1_impl_0_out);

   Delay1No358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_0_out,
                 Y => Delay1No358_out);

SharedReg394_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg395_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg395_out;
SharedReg392_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg392_out;
SharedReg398_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg398_out;
   MUX_Product26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg395_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg392_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg398_out_to_MUX_Product26_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product26_1_impl_1_out);

   Delay1No359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_1_impl_1_out,
                 Y => Delay1No359_out);

Delay1No360_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast <= Delay1No360_out;
Delay1No361_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast <= Delay1No361_out;
   Product26_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product26_2_impl_out,
                 X => Delay1No360_out_to_Product26_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No361_out_to_Product26_2_impl_parent_implementedSystem_port_1_cast);

SharedReg28_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg28_out;
SharedReg363_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg363_out;
SharedReg263_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg321_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg321_out;
   MUX_Product26_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg28_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg363_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg263_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg321_out_to_MUX_Product26_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product26_2_impl_0_out);

   Delay1No360_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_2_impl_0_out,
                 Y => Delay1No360_out);

SharedReg388_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg398_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg398_out;
SharedReg394_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg394_out;
SharedReg400_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
   MUX_Product26_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg398_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg394_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Product26_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product26_2_impl_1_out);

   Delay1No361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product26_2_impl_1_out,
                 Y => Delay1No361_out);

Delay1No362_out_to_Product27_0_impl_parent_implementedSystem_port_0_cast <= Delay1No362_out;
Delay1No363_out_to_Product27_0_impl_parent_implementedSystem_port_1_cast <= Delay1No363_out;
   Product27_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product27_0_impl_out,
                 X => Delay1No362_out_to_Product27_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No363_out_to_Product27_0_impl_parent_implementedSystem_port_1_cast);

SharedReg323_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg323_out;
SharedReg28_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg324_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg324_out;
SharedReg343_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg343_out;
   MUX_Product27_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg323_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg324_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Product27_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_0_impl_0_out);

   Delay1No362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_0_impl_0_out,
                 Y => Delay1No362_out);

SharedReg400_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg400_out;
SharedReg388_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg393_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg393_out;
SharedReg105_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product27_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg393_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product27_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_0_impl_1_out);

   Delay1No363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_0_impl_1_out,
                 Y => Delay1No363_out);

Delay1No364_out_to_Product27_1_impl_parent_implementedSystem_port_0_cast <= Delay1No364_out;
Delay1No365_out_to_Product27_1_impl_parent_implementedSystem_port_1_cast <= Delay1No365_out;
   Product27_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product27_1_impl_out,
                 X => Delay1No364_out_to_Product27_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No365_out_to_Product27_1_impl_parent_implementedSystem_port_1_cast);

SharedReg160_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg160_out;
SharedReg383_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg383_out;
SharedReg28_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg327_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg327_out;
   MUX_Product27_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg160_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg383_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg28_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg327_out_to_MUX_Product27_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_1_impl_0_out);

   Delay1No364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_1_impl_0_out,
                 Y => Delay1No364_out);

SharedReg169_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg397_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg397_out;
SharedReg388_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg388_out;
SharedReg393_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg393_out;
   MUX_Product27_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg397_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg388_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg393_out_to_MUX_Product27_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_1_impl_1_out);

   Delay1No365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_1_impl_1_out,
                 Y => Delay1No365_out);

Delay1No366_out_to_Product27_2_impl_parent_implementedSystem_port_0_cast <= Delay1No366_out;
Delay1No367_out_to_Product27_2_impl_parent_implementedSystem_port_1_cast <= Delay1No367_out;
   Product27_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product27_2_impl_out,
                 X => Delay1No366_out_to_Product27_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No367_out_to_Product27_2_impl_parent_implementedSystem_port_1_cast);

SharedReg29_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg29_out;
SharedReg322_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg322_out;
SharedReg348_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg348_out;
SharedReg363_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg363_out;
   MUX_Product27_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg29_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg322_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg348_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg363_out_to_MUX_Product27_2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_2_impl_0_out);

   Delay1No366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_2_impl_0_out,
                 Y => Delay1No366_out);

SharedReg388_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg393_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg393_out;
SharedReg351_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg351_out;
SharedReg400_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
   MUX_Product27_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg393_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg351_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Product27_2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_2_impl_1_out);

   Delay1No367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_2_impl_1_out,
                 Y => Delay1No367_out);

Delay1No368_out_to_Product48_0_impl_parent_implementedSystem_port_0_cast <= Delay1No368_out;
Delay1No369_out_to_Product48_0_impl_parent_implementedSystem_port_1_cast <= Delay1No369_out;
   Product48_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product48_0_impl_out,
                 X => Delay1No368_out_to_Product48_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No369_out_to_Product48_0_impl_parent_implementedSystem_port_1_cast);

SharedReg365_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg365_out;
SharedReg29_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg3_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg114_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg114_out;
   MUX_Product48_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg365_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg3_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg114_out_to_MUX_Product48_0_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product48_0_impl_0_out);

   Delay1No368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_0_impl_0_out,
                 Y => Delay1No368_out);

SharedReg400_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg400_out;
SharedReg388_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg388_out;
SharedReg113_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg113_out;
SharedReg105_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Product48_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg388_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg113_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Product48_0_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product48_0_impl_1_out);

   Delay1No369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_0_impl_1_out,
                 Y => Delay1No369_out);

Delay1No370_out_to_Product48_1_impl_parent_implementedSystem_port_0_cast <= Delay1No370_out;
Delay1No371_out_to_Product48_1_impl_parent_implementedSystem_port_1_cast <= Delay1No371_out;
   Product48_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product48_1_impl_out,
                 X => Delay1No370_out_to_Product48_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No371_out_to_Product48_1_impl_parent_implementedSystem_port_1_cast);

SharedReg111_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg356_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg356_out;
SharedReg29_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg3_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg3_out;
   MUX_Product48_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg356_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg29_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg3_out_to_MUX_Product48_1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product48_1_impl_0_out);

   Delay1No370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_1_impl_0_out,
                 Y => Delay1No370_out);

SharedReg169_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg169_out;
SharedReg400_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg400_out;
SharedReg388_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg388_out;
SharedReg110_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg110_out;
   MUX_Product48_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg169_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg400_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg388_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Product48_1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product48_1_impl_1_out);

   Delay1No371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_1_impl_1_out,
                 Y => Delay1No371_out);

Delay1No372_out_to_Product48_2_impl_parent_implementedSystem_port_0_cast <= Delay1No372_out;
Delay1No373_out_to_Product48_2_impl_parent_implementedSystem_port_1_cast <= Delay1No373_out;
   Product48_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product48_2_impl_out,
                 X => Delay1No372_out_to_Product48_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No373_out_to_Product48_2_impl_parent_implementedSystem_port_1_cast);

SharedReg3_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg3_out;
SharedReg30_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg30_out;
SharedReg386_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg386_out;
   MUX_Product48_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg3_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg386_out_to_MUX_Product48_2_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product48_2_impl_0_LUT_out,
                 oMux => MUX_Product48_2_impl_0_out);

   Delay1No372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_2_impl_0_out,
                 Y => Delay1No372_out);

SharedReg351_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg351_out;
SharedReg385_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg385_out;
SharedReg388_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg388_out;
   MUX_Product48_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg351_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg385_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg388_out_to_MUX_Product48_2_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product48_2_impl_1_LUT_out,
                 oMux => MUX_Product48_2_impl_1_out);

   Delay1No373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product48_2_impl_1_out,
                 Y => Delay1No373_out);

Delay1No374_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No374_out;
Delay1No375_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No375_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No374_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No375_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

   Delay1No374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => Delay1No374_out);

   Delay1No375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => Delay1No375_out);
   Constant_0_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);

   Delay111No1_instance: Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=107 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => Delay111No1_out);

   Delay114No_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => Delay114No_out);

   Delay114No1_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => Delay114No1_out);

   Delay114No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => Delay114No2_out);

   Delay112No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => Delay112No2_out);

   Delay113No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay113No1_out);

   Delay111No3_instance: Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=108 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => Delay111No3_out);

   Delay2No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => Delay2No1_out);

   Delay100No1_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => Delay100No1_out);

   Delay5No9_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => Delay5No9_out);

   Delay103No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => Delay103No_out);

   Delay103No1_instance: Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=102 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => Delay103No1_out);

   Delay103No2_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => Delay103No2_out);

   Delay114No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => Delay114No3_out);

   Delay114No4_instance: Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=107 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => Delay114No4_out);

   Delay114No5_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => Delay114No5_out);

   Delay115No_instance: Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=111 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => Delay115No_out);

   Delay115No1_instance: Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=111 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => Delay115No1_out);

   Delay115No2_instance: Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=111 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => Delay115No2_out);

   Delay115No3_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => Delay115No3_out);

   Delay115No4_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => Delay115No4_out);

   Delay115No5_instance: Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=111 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => Delay115No5_out);

   Delay110No_instance: Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=103 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => Delay110No_out);

   Delay110No2_instance: Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=105 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => Delay110No2_out);

   Delay3No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay3No6_out);

   Delay3No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => Delay3No7_out);

   Delay3No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => Delay3No8_out);

   Delay14No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => Delay14No_out);

   Delay14No2_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => Delay14No2_out);

   Delay7No54_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => Delay7No54_out);

   Delay7No55_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => Delay7No55_out);

   Delay14No5_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => Delay14No5_out);

   Delay20No_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay20No_out);

   Delay20No1_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay20No1_out);

   Delay20No2_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay20No2_out);

   Delay6No5_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay6No5_out);

   Delay3No9_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => Delay3No9_out);

   Delay3No10_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay3No10_out);

   Delay6No6_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => Delay6No6_out);

   Delay6No7_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => Delay6No7_out);

   Delay6No8_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay6No8_out);

   Delay2No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => Delay2No9_out);

   Delay2No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => Delay2No10_out);

   Delay2No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => Delay2No11_out);

   Delay2No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => Delay2No12_out);

   Delay2No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => Delay2No13_out);

   Delay2No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay2No14_out);

   Delay11No_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => Delay11No_out);

   Delay11No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => Delay11No1_out);

   Delay7No58_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => Delay7No58_out);

   Delay16No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => Delay16No_out);

   Delay16No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => Delay16No1_out);

   Delay11No8_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => Delay11No8_out);

   Delay5No13_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => Delay5No13_out);

   Delay5No14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => Delay5No14_out);

   Delay3No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => Delay3No15_out);

   Delay3No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => Delay3No16_out);

   Delay6No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => Delay6No18_out);

   Delay6No19_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => Delay6No19_out);

   Delay6No20_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => Delay6No20_out);

   Delay3No21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => Delay3No21_out);

   Delay3No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => Delay3No24_out);

   Delay3No25_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => Delay3No25_out);

   Delay10No21_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay10No21_out);

   Delay10No22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => Delay10No22_out);

   Delay8No21_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => Delay8No21_out);

   Delay8No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => Delay8No22_out);

   Delay2No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => Delay2No41_out);

   Delay7No60_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => Delay7No60_out);

   Delay2No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => Delay2No43_out);

   Delay2No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => Delay2No44_out);

   Delay8No24_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => Delay8No24_out);

   Delay8No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => Delay8No26_out);

   Delay8No27_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => Delay8No27_out);

   Delay8No28_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => Delay8No28_out);

   Delay5No18_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => Delay5No18_out);

   Delay5No19_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => Delay5No19_out);

   Delay5No23_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => Delay5No23_out);

   Delay15No_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => Delay15No_out);

   Delay15No1_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => Delay15No1_out);

   Delay11No9_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => Delay11No9_out);

   Delay11No10_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => Delay11No10_out);

   Delay11No11_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => Delay11No11_out);

   Delay2No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => Delay2No45_out);

   Delay21No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => Delay21No1_out);

   Delay18No2_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => Delay18No2_out);

   Delay22No_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => Delay22No_out);

   Delay22No1_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay22No1_out);

   Delay22No2_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => Delay22No2_out);

   Delay17No_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => Delay17No_out);

   Delay17No1_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => Delay17No1_out);

   Delay17No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => Delay17No2_out);

   Delay12No18_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => Delay12No18_out);

   Delay12No19_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => Delay12No19_out);

   Delay12No20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => Delay12No20_out);

   Delay17No3_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => Delay17No3_out);

   Delay17No5_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => Delay17No5_out);

   Delay12No25_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => Delay12No25_out);

   Delay18No3_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => Delay18No3_out);

   Delay18No4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => Delay18No4_out);

   Delay18No5_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => Delay18No5_out);

   Delay3No27_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => Delay3No27_out);

   Delay3No30_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => Delay3No30_out);

   Delay3No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => Delay3No31_out);

   Delay3No32_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => Delay3No32_out);

   Delay4No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => Delay4No7_out);

   Delay4No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => Delay4No8_out);

   Delay2No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => Delay2No54_out);

   Delay2No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => Delay2No56_out);

   Delay73No_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => Delay73No_out);

   Delay73No1_instance: Delay_34_DelayLength_72_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=72 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => Delay73No1_out);

   Delay73No2_instance: Delay_34_DelayLength_59_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=59 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => Delay73No2_out);

   Delay68No_instance: Delay_34_DelayLength_54_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=54 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => Delay68No_out);

   Delay68No1_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => Delay68No1_out);

   Delay71No_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => Delay71No_out);

   Delay71No1_instance: Delay_34_DelayLength_69_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=69 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => Delay71No1_out);

   Delay71No2_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => Delay71No2_out);

   Delay95No_instance: Delay_34_DelayLength_91_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=91 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => Delay95No_out);

   Delay95No1_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => Delay95No1_out);

   Delay95No2_instance: Delay_34_DelayLength_80_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=80 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => Delay95No2_out);

   Delay57No_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => Delay57No_out);

   Delay57No2_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => Delay57No2_out);

   Delay51No_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay51No_out);

   Delay51No1_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => Delay51No1_out);

   Delay51No2_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => Delay51No2_out);

   Delay3No33_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => Delay3No33_out);

   Delay3No34_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => Delay3No34_out);

   Delay36No_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => Delay36No_out);

   Delay36No1_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => Delay36No1_out);

   Delay37No_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => Delay37No_out);

   Delay37No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => Delay37No1_out);

   Delay37No2_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => Delay37No2_out);

   Delay32No_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => Delay32No_out);

   Delay32No1_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => Delay32No1_out);

   Delay32No2_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => Delay32No2_out);

   Delay27No_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => Delay27No_out);

   Delay27No1_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => Delay27No1_out);

   Delay27No2_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => Delay27No2_out);

   Delay4No46_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => Delay4No46_out);

   Delay4No49_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => Delay4No49_out);

   Delay2No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => Delay2No63_out);

   Delay2No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => Delay2No65_out);

   Delay87No_instance: Delay_34_DelayLength_76_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=76 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => Delay87No_out);

   Delay87No1_instance: Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=85 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => Delay87No1_out);

   Delay87No2_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => Delay87No2_out);

   Delay11No13_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => Delay11No13_out);

   Delay11No14_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => Delay11No14_out);

   Delay90No_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => Delay90No_out);

   Delay90No1_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => Delay90No1_out);

   Delay90No2_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => Delay90No2_out);

   MUX_Inv_11_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_11_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_11_0_0_LUT_out);

   MUX_Inv_12_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_12_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_12_0_0_LUT_out);

   MUX_Inv_13_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_13_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_13_0_0_LUT_out);

   MUX_Inv_21_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_21_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_21_0_0_LUT_out);

   MUX_Inv_22_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_22_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_22_0_0_LUT_out);

   MUX_Inv_23_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_23_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_23_0_0_LUT_out);

   MUX_Inv_31_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_31_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_31_0_0_LUT_out);

   MUX_Inv_32_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_32_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_32_0_0_LUT_out);

   MUX_Inv_33_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_33_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_33_0_0_LUT_out);

   MUX_Inv_41_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_41_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_41_0_0_LUT_out);

   MUX_Inv_42_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_42_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_42_0_0_LUT_out);

   MUX_Inv_43_0_0_LUT_instance: GenericLut_LUTData_MUX_Inv_43_0_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Inv_43_0_0_LUT_out);

   MUX_Subtract5_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract5_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract5_2_impl_0_LUT_out);

   MUX_Subtract5_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract5_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract5_2_impl_1_LUT_out);

   MUX_Add9_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add9_2_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add9_2_impl_0_LUT_out);

   MUX_Add9_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add9_2_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add9_2_impl_1_LUT_out);

   MUX_Divide_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Divide_0_impl_0_LUT_out);

   MUX_Divide_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Divide_0_impl_1_LUT_out);

   MUX_Product48_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product48_2_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product48_2_impl_0_LUT_out);

   MUX_Product48_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product48_2_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product48_2_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_0_impl_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_1_impl_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_2_impl_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_0_impl_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_1_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_2_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_0_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_1_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_2_impl_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_0_impl_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_1_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_2_impl_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_0_impl_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_1_impl_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_2_impl_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_0_impl_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_1_impl_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_2_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_0_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_1_impl_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_2_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_0_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_1_impl_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_2_impl_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_0_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_1_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_2_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_0_impl_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_1_impl_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_2_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_0_impl_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_1_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_2_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_0_impl_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_1_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_2_impl_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_0_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_110_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=110 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_1_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_2_impl_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_1_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_2_impl_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=108 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_2_impl_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_1_impl_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_108_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=108 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_2_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_110_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=110 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_0_impl_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_1_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add131_0_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_111_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=111 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add131_1_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_105_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=105 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_0_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_1_impl_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_2_impl_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add210_0_impl_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add210_1_impl_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add20_2_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_89_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=89 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add21_0_impl_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=92 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add21_1_impl_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_92_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=92 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_0_impl_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_1_impl_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_2_impl_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add25_0_impl_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add25_1_impl_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add25_2_impl_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add28_0_impl_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add28_1_impl_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add28_2_impl_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add71_2_impl_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add81_0_impl_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add81_1_impl_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product112_1_impl_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_0_impl_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_1_impl_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product113_2_impl_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_0_impl_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_1_impl_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product102_2_impl_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_0_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_1_impl_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_2_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product131_0_impl_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product131_1_impl_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product131_2_impl_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product371_2_impl_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product381_0_impl_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product381_1_impl_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product391_2_impl_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product411_0_impl_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product411_2_impl_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product421_0_impl_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product421_1_impl_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product421_2_impl_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product441_0_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product441_1_impl_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product441_2_impl_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product461_0_impl_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product461_1_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product461_2_impl_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product481_0_impl_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product481_1_impl_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product481_2_impl_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product511_0_impl_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product511_1_impl_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product511_2_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product521_0_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product521_1_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product521_2_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_0_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_1_impl_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_2_impl_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product57_0_impl_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product57_1_impl_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product57_2_impl_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product59_0_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product59_1_impl_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product59_2_impl_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product61_0_impl_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product61_1_impl_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product61_2_impl_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product62_0_impl_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product62_1_impl_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product62_2_impl_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product63_0_impl_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product63_1_impl_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product63_2_impl_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product64_0_impl_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product64_1_impl_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product64_2_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product66_0_impl_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product66_1_impl_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product66_2_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product67_0_impl_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product67_1_impl_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product67_2_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product68_0_impl_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product68_1_impl_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product68_2_impl_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product711_0_impl_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product711_1_impl_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product711_2_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product70_0_impl_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product70_1_impl_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product70_2_impl_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product71_0_impl_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product71_1_impl_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product71_2_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product76_0_impl_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product76_1_impl_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product76_2_impl_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product911_0_impl_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product911_1_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product911_2_impl_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_0_impl_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_1_impl_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_2_impl_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract1_2_impl_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract11_1_impl_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_0_impl_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_1_impl_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_2_impl_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract5_2_impl_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add32_0_impl_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add32_2_impl_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add211_2_impl_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add6_2_impl_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_2_impl_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_123_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=123 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_0_impl_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_0_impl_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_1_impl_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_2_impl_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product14_0_impl_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product14_1_impl_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product14_2_impl_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=67 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_0_impl_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_1_impl_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product26_2_impl_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product27_0_impl_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product27_1_impl_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product27_2_impl_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product48_0_impl_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product48_1_impl_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product48_2_impl_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => SharedReg400_out);
end architecture;

