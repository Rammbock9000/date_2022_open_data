--------------------------------------------------------------------------------
--                         ModuloCounter_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_4_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of ModuloCounter_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(1 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 3 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2400610_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2400612)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2400610_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2400610_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2400615
--                  (IntAdderAlternative_27_f250_uid2400619)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2400615 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2400615 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2400622
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2400622 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2400622 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2400625
--                   (IntAdderClassical_34_f250_uid2400627)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2400625 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2400625 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2400610
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2400610 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2400610 is
   component FPAdd_8_23_uid2400610_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2400615 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2400622 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2400625 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2400610_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2400615  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2400622  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2400625  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2400610 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2400610  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_4_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
         iS_3 when "11",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2401370
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2401370 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2401370 is
signal XX_m2401371 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2401371 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2401371 <= X ;
   YY_m2401371 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2401374
--                   (IntAdderClassical_33_f500_uid2401376)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2401374 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2401374 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2401370 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2401374 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2401370  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2401374  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2401457_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2401459)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2401457_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2401457_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2401462
--                  (IntAdderAlternative_27_f250_uid2401466)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2401462 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2401462 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2401469
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2401469 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2401469 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2401472
--                   (IntAdderClassical_34_f250_uid2401474)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2401472 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2401472 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2401457
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2401457 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2401457 is
   component FPAdd_8_23_uid2401457_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2401462 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2401469 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2401472 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2401457_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2401462  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2401469  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2401472  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2401457 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2401457  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_3_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_3_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(1 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_3_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00",
         iS_1 when "01",
         iS_2 when "10",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_2_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(0 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0",
         iS_1 when "1",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--            GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "1" when "00",
      "0" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--   GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "10" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "10" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "10" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "00" when "01",
      "01" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "00" when "01",
      "01" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "10" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "01" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "00" when "01",
      "00" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "01" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "00" when "01",
      "00" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "01" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "01" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "01" when "00",
      "00" when "01",
      "00" when "10",
      "10" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "00" when "00",
      "00" when "01",
      "10" when "10",
      "01" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "0" when "10",
      "1" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "0" when "10",
      "1" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "0" when "10",
      "1" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "0" when "01",
      "0" when "10",
      "1" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "00" when "01",
      "01" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "00" when "01",
      "01" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "01" when "01",
      "00" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(1 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "10" when "00",
      "01" when "01",
      "00" when "10",
      "00" when "11",
      "00" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(1 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          o0 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1 is
signal t_in : std_logic_vector(1 downto 0) := (others => '0');
signal t_out : std_logic_vector(0 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   with t_in select t_out <= 
      "0" when "00",
      "1" when "01",
      "0" when "10",
      "0" when "11",
      "0" when others;

   o0 <= t_out(0);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(1 downto 0);
          Output : out std_logic_vector(0 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
   component GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             o0 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
   instLUT: GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 o0 => Output0_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re : in std_logic_vector(31 downto 0);
          x0_im : in std_logic_vector(31 downto 0);
          x1_re : in std_logic_vector(31 downto 0);
          x1_im : in std_logic_vector(31 downto 0);
          x2_re : in std_logic_vector(31 downto 0);
          x2_im : in std_logic_vector(31 downto 0);
          x3_re : in std_logic_vector(31 downto 0);
          x3_im : in std_logic_vector(31 downto 0);
          x4_re : in std_logic_vector(31 downto 0);
          x4_im : in std_logic_vector(31 downto 0);
          x5_re : in std_logic_vector(31 downto 0);
          x5_im : in std_logic_vector(31 downto 0);
          x6_re : in std_logic_vector(31 downto 0);
          x6_im : in std_logic_vector(31 downto 0);
          x7_re : in std_logic_vector(31 downto 0);
          x7_im : in std_logic_vector(31 downto 0);
          x8_re : in std_logic_vector(31 downto 0);
          x8_im : in std_logic_vector(31 downto 0);
          x9_re : in std_logic_vector(31 downto 0);
          x9_im : in std_logic_vector(31 downto 0);
          x10_re : in std_logic_vector(31 downto 0);
          x10_im : in std_logic_vector(31 downto 0);
          x11_re : in std_logic_vector(31 downto 0);
          x11_im : in std_logic_vector(31 downto 0);
          x12_re : in std_logic_vector(31 downto 0);
          x12_im : in std_logic_vector(31 downto 0);
          x13_re : in std_logic_vector(31 downto 0);
          x13_im : in std_logic_vector(31 downto 0);
          x14_re : in std_logic_vector(31 downto 0);
          x14_im : in std_logic_vector(31 downto 0);
          x15_re : in std_logic_vector(31 downto 0);
          x15_im : in std_logic_vector(31 downto 0);
          y0_re : out std_logic_vector(31 downto 0);
          y0_im : out std_logic_vector(31 downto 0);
          y1_re : out std_logic_vector(31 downto 0);
          y1_im : out std_logic_vector(31 downto 0);
          y2_re : out std_logic_vector(31 downto 0);
          y2_im : out std_logic_vector(31 downto 0);
          y3_re : out std_logic_vector(31 downto 0);
          y3_im : out std_logic_vector(31 downto 0);
          y4_re : out std_logic_vector(31 downto 0);
          y4_im : out std_logic_vector(31 downto 0);
          y5_re : out std_logic_vector(31 downto 0);
          y5_im : out std_logic_vector(31 downto 0);
          y6_re : out std_logic_vector(31 downto 0);
          y6_im : out std_logic_vector(31 downto 0);
          y7_re : out std_logic_vector(31 downto 0);
          y7_im : out std_logic_vector(31 downto 0);
          y8_re : out std_logic_vector(31 downto 0);
          y8_im : out std_logic_vector(31 downto 0);
          y9_re : out std_logic_vector(31 downto 0);
          y9_im : out std_logic_vector(31 downto 0);
          y10_re : out std_logic_vector(31 downto 0);
          y10_im : out std_logic_vector(31 downto 0);
          y11_re : out std_logic_vector(31 downto 0);
          y11_im : out std_logic_vector(31 downto 0);
          y12_re : out std_logic_vector(31 downto 0);
          y12_im : out std_logic_vector(31 downto 0);
          y13_re : out std_logic_vector(31 downto 0);
          y13_im : out std_logic_vector(31 downto 0);
          y14_re : out std_logic_vector(31 downto 0);
          y14_im : out std_logic_vector(31 downto 0);
          y15_re : out std_logic_vector(31 downto 0);
          y15_im : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_4_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(1 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_4_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_3_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(1 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_2_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(0 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(1 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(1 downto 0);
             Output : out std_logic_vector(0 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount41_out : std_logic_vector(1 downto 0) := (others => '0');
signal x0_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add15_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add16_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add22_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add112_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add112_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add121_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add33_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add34_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add34_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add124_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add124_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add124_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add37_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add37_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add127_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add129_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add129_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add130_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add130_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add42_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add42_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add42_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product13_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product7_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product17_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product27_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract8_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract10_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product30_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product30_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract11_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add53_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add53_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add54_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product42_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product42_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product114_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product313_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product313_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract14_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract14_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add57_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add57_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add58_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add58_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add58_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add59_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add59_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add59_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product118_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product118_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product118_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product217_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product217_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product217_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product317_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product317_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product317_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract19_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract19_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product219_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product219_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product219_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product49_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product49_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product220_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract21_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product122_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product122_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product221_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product221_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product321_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product321_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract22_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product223_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product223_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product223_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract24_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product53_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product53_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product125_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product125_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product125_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product324_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product324_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract25_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract25_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add67_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add67_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add67_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add68_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product127_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract36_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract36_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract36_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product237_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product237_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product237_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product337_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product337_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product337_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product67_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product67_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product338_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product338_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product338_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product68_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product68_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product339_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product339_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product339_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product145_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product145_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product145_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product244_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product244_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product244_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract46_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract47_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product148_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product148_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product148_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product347_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product347_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product347_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract50_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract50_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract111_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract111_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract116_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract116_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract57_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract117_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract61_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract61_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract61_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract121_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract121_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract125_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract125_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract125_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract66_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract66_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract66_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract126_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract126_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract126_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract135_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract135_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract135_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract137_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract137_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract137_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract79_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract79_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract79_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract139_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract139_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract139_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant12_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant10_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant19_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant20_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant110_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant21_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant111_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant22_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant112_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant23_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant113_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant24_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant114_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant25_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant115_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant26_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant116_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant27_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant117_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant28_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant118_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant29_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant119_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant30_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant120_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant31_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant121_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant32_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant122_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant33_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant123_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant34_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant124_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant35_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant125_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant36_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant126_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant37_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant127_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant38_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant128_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant39_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant129_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant40_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant130_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant41_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant131_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant42_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant132_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant43_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant133_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant44_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant134_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant45_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant135_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant46_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant136_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant47_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant137_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant48_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant138_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant49_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant139_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant50_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant140_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant51_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant141_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant52_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant142_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant53_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant143_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant54_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant144_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant55_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant145_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant56_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant146_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant57_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant147_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add57_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add57_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add58_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add58_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add59_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add59_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Add67_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Add67_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product237_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product237_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product337_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product337_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product67_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product67_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product338_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product338_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product68_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product68_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product339_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product339_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product145_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product145_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product244_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product244_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Product148_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product148_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product347_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Product347_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract126_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract126_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract135_impl_0_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract135_impl_1_LUT_out : std_logic_vector(1 downto 0) := (others => '0');
signal MUX_Subtract137_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract137_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract79_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract79_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract139_impl_0_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal MUX_Subtract139_impl_1_LUT_out : std_logic_vector(0 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y1_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y1_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y2_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y2_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y3_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y3_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y4_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y4_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y5_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y5_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y6_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y6_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y7_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y7_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y8_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y8_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y9_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y9_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y10_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y10_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y11_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y11_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y12_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y12_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y13_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y13_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y14_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y14_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y15_re_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y15_im_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No63_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No57_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No66_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No1_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add15_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add15_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add16_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add16_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add9_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add9_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add18_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add18_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No4_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No13_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add22_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add22_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add112_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add112_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add121_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add121_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add33_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add33_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add34_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add34_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No43_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add124_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add124_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add37_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add37_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No60_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add127_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add127_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No56_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No48_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add129_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add129_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add40_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add40_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No3_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No52_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add130_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add130_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add42_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add42_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No54_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No1_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No2_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No2_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No76_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No3_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product31_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product31_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No39_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product6_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product6_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product13_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product13_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product23_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product23_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product33_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product33_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product7_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product7_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product10_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product10_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product17_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product17_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product27_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product27_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No14_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No24_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product37_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product37_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No14_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No15_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No27_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Subtract8_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Subtract8_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No1_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Subtract10_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Subtract10_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No44_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product30_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product30_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product210_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product210_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product310_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product310_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Add53_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Add53_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Add54_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Add54_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product42_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product42_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product114_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product114_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product213_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product213_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product313_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product313_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Subtract14_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Subtract14_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Add57_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Add57_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Add58_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Add58_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No67_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Add59_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Add59_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product118_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product118_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No6_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product217_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product217_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product317_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product317_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Subtract19_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Subtract19_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No2_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No49_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product219_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product219_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No9_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No50_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product49_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product49_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay21No31_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No9_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No10_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product220_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product220_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Subtract21_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Subtract21_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No51_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product122_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product122_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product221_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product221_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product321_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product321_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Subtract22_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Subtract22_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No68_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product223_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product223_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay22No_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No8_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Subtract24_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Subtract24_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No53_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No55_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product53_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product53_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product125_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product125_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product324_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product324_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Subtract25_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Subtract25_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Add67_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Add67_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Add68_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Add68_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Product55_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Product55_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product127_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product127_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Product226_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Product226_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product326_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product326_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Subtract36_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Subtract36_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Product237_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Product237_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Product337_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Product337_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product67_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product67_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No34_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No72_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product338_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product338_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No73_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No35_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product68_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product68_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No32_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No17_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No74_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product339_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product339_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No75_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay7No18_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay36No33_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product145_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product145_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No3_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No29_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Product244_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Product244_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay8No4_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Subtract46_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Subtract46_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Subtract47_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Subtract47_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Product148_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Product148_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product148_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product148_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product148_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product148_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Product347_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Product347_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product347_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product347_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product347_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product347_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Subtract50_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Subtract50_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No9_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Subtract111_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Subtract111_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No36_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Subtract116_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Subtract116_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No40_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Subtract57_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Subtract57_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Subtract117_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Subtract117_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No58_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Subtract61_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Subtract61_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Subtract121_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Subtract121_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Subtract125_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Subtract125_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Subtract66_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Subtract66_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Subtract126_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Subtract126_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Subtract135_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Subtract135_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No3_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No12_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Subtract137_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Subtract137_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract137_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract137_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract137_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract137_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Subtract79_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Subtract79_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No7_out_to_MUX_Subtract79_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Subtract79_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No16_out_to_MUX_Subtract79_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Subtract79_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Subtract139_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Subtract139_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No8_out_to_MUX_Subtract139_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Subtract139_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay2No17_out_to_MUX_Subtract139_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Subtract139_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount41_instance: ModuloCounter_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount41_out);
x0_re_IEEE <= x0_re;
   x0_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_out,
                 X => x0_re_IEEE);
x0_im_IEEE <= x0_im;
   x0_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_out,
                 X => x0_im_IEEE);
x1_re_IEEE <= x1_re;
   x1_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_out,
                 X => x1_re_IEEE);
x1_im_IEEE <= x1_im;
   x1_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_out,
                 X => x1_im_IEEE);
x2_re_IEEE <= x2_re;
   x2_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_out,
                 X => x2_re_IEEE);
x2_im_IEEE <= x2_im;
   x2_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_out,
                 X => x2_im_IEEE);
x3_re_IEEE <= x3_re;
   x3_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_out,
                 X => x3_re_IEEE);
x3_im_IEEE <= x3_im;
   x3_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_out,
                 X => x3_im_IEEE);
x4_re_IEEE <= x4_re;
   x4_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_out,
                 X => x4_re_IEEE);
x4_im_IEEE <= x4_im;
   x4_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_out,
                 X => x4_im_IEEE);
x5_re_IEEE <= x5_re;
   x5_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_out,
                 X => x5_re_IEEE);
x5_im_IEEE <= x5_im;
   x5_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_out,
                 X => x5_im_IEEE);
x6_re_IEEE <= x6_re;
   x6_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_out,
                 X => x6_re_IEEE);
x6_im_IEEE <= x6_im;
   x6_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_out,
                 X => x6_im_IEEE);
x7_re_IEEE <= x7_re;
   x7_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_out,
                 X => x7_re_IEEE);
x7_im_IEEE <= x7_im;
   x7_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_out,
                 X => x7_im_IEEE);
x8_re_IEEE <= x8_re;
   x8_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_out,
                 X => x8_re_IEEE);
x8_im_IEEE <= x8_im;
   x8_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_out,
                 X => x8_im_IEEE);
x9_re_IEEE <= x9_re;
   x9_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_out,
                 X => x9_re_IEEE);
x9_im_IEEE <= x9_im;
   x9_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_out,
                 X => x9_im_IEEE);
x10_re_IEEE <= x10_re;
   x10_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_out,
                 X => x10_re_IEEE);
x10_im_IEEE <= x10_im;
   x10_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_out,
                 X => x10_im_IEEE);
x11_re_IEEE <= x11_re;
   x11_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_out,
                 X => x11_re_IEEE);
x11_im_IEEE <= x11_im;
   x11_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_out,
                 X => x11_im_IEEE);
x12_re_IEEE <= x12_re;
   x12_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_out,
                 X => x12_re_IEEE);
x12_im_IEEE <= x12_im;
   x12_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_out,
                 X => x12_im_IEEE);
x13_re_IEEE <= x13_re;
   x13_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_out,
                 X => x13_re_IEEE);
x13_im_IEEE <= x13_im;
   x13_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_out,
                 X => x13_im_IEEE);
x14_re_IEEE <= x14_re;
   x14_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_out,
                 X => x14_re_IEEE);
x14_im_IEEE <= x14_im;
   x14_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_out,
                 X => x14_im_IEEE);
x15_re_IEEE <= x15_re;
   x15_re_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_out,
                 X => x15_re_IEEE);
x15_im_IEEE <= x15_im;
   x15_im_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_out,
                 X => x15_im_IEEE);
   y0_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_IEEE,
                 X => Delay1No_out);
y0_re <= y0_re_IEEE;

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => Delay1No_out);
   y0_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_IEEE,
                 X => Delay1No1_out);
y0_im <= y0_im_IEEE;

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => Delay1No1_out);
   y1_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_IEEE,
                 X => Delay1No2_out);
y1_re <= y1_re_IEEE;

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => Delay1No2_out);
   y1_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_IEEE,
                 X => Delay1No3_out);
y1_im <= y1_im_IEEE;

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay1No3_out);
   y2_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_IEEE,
                 X => Delay1No4_out);
y2_re <= y2_re_IEEE;

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => Delay1No4_out);
   y2_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_IEEE,
                 X => Delay1No5_out);
y2_im <= y2_im_IEEE;

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay1No5_out);
   y3_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_IEEE,
                 X => Delay1No6_out);
y3_re <= y3_re_IEEE;

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No6_out);
   y3_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_IEEE,
                 X => Delay1No7_out);
y3_im <= y3_im_IEEE;

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay1No7_out);
   y4_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_IEEE,
                 X => Delay1No8_out);
y4_re <= y4_re_IEEE;

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => Delay1No8_out);
   y4_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_IEEE,
                 X => Delay1No9_out);
y4_im <= y4_im_IEEE;

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay1No9_out);
   y5_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_IEEE,
                 X => Delay1No10_out);
y5_re <= y5_re_IEEE;

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay1No10_out);
   y5_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_IEEE,
                 X => Delay1No11_out);
y5_im <= y5_im_IEEE;

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => Delay1No11_out);
   y6_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_IEEE,
                 X => Delay1No12_out);
y6_re <= y6_re_IEEE;

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => Delay1No12_out);
   y6_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_IEEE,
                 X => Delay1No13_out);
y6_im <= y6_im_IEEE;

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => Delay1No13_out);
   y7_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_IEEE,
                 X => Delay1No14_out);
y7_re <= y7_re_IEEE;

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => Delay1No14_out);
   y7_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_IEEE,
                 X => Delay1No15_out);
y7_im <= y7_im_IEEE;

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => Delay1No15_out);
   y8_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_IEEE,
                 X => Delay1No16_out);
y8_re <= y8_re_IEEE;

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => Delay1No16_out);
   y8_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_IEEE,
                 X => Delay1No17_out);
y8_im <= y8_im_IEEE;

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => Delay1No17_out);
   y9_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_IEEE,
                 X => Delay1No18_out);
y9_re <= y9_re_IEEE;

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => Delay1No18_out);
   y9_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_IEEE,
                 X => Delay1No19_out);
y9_im <= y9_im_IEEE;

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => Delay1No19_out);
   y10_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_IEEE,
                 X => Delay1No20_out);
y10_re <= y10_re_IEEE;

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => Delay1No20_out);
   y10_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_IEEE,
                 X => Delay1No21_out);
y10_im <= y10_im_IEEE;

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => Delay1No21_out);
   y11_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_IEEE,
                 X => Delay1No22_out);
y11_re <= y11_re_IEEE;

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => Delay1No22_out);
   y11_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_IEEE,
                 X => Delay1No23_out);
y11_im <= y11_im_IEEE;

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => Delay1No23_out);
   y12_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_IEEE,
                 X => Delay1No24_out);
y12_re <= y12_re_IEEE;

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => Delay1No24_out);
   y12_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_IEEE,
                 X => Delay1No25_out);
y12_im <= y12_im_IEEE;

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => Delay1No25_out);
   y13_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_IEEE,
                 X => Delay1No26_out);
y13_re <= y13_re_IEEE;

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => Delay1No26_out);
   y13_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_IEEE,
                 X => Delay1No27_out);
y13_im <= y13_im_IEEE;

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => Delay1No27_out);
   y14_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_IEEE,
                 X => Delay1No28_out);
y14_re <= y14_re_IEEE;

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => Delay1No28_out);
   y14_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_IEEE,
                 X => Delay1No29_out);
y14_im <= y14_im_IEEE;

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => Delay1No29_out);
   y15_re_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_IEEE,
                 X => Delay1No30_out);
y15_re <= y15_re_IEEE;

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => Delay1No30_out);
   y15_im_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_IEEE,
                 X => Delay1No31_out);
y15_im <= y15_im_IEEE;

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_impl_out,
                 X => Delay1No32_out_to_Add2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_impl_parent_implementedSystem_port_1_cast);

SharedReg54_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg54_out;
SharedReg_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg3_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg48_out;
   MUX_Add2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg54_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg3_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg48_out_to_MUX_Add2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add2_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_impl_0_out,
                 Y => Delay1No32_out);

Delay2No63_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast <= Delay2No63_out;
SharedReg16_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg19_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg50_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg50_out;
   MUX_Add2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No63_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg19_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg50_out_to_MUX_Add2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add2_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add11_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add11_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add11_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_impl_out,
                 X => Delay1No34_out_to_Add11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add11_impl_parent_implementedSystem_port_1_cast);

Delay2No57_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_1_cast <= Delay2No57_out;
SharedReg1_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg88_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
Delay3No_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_4_cast <= Delay3No_out;
   MUX_Add11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No57_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No_out_to_MUX_Add11_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add11_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_impl_0_out,
                 Y => Delay1No34_out);

Delay2No66_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_1_cast <= Delay2No66_out;
SharedReg17_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg108_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_3_cast <= SharedReg108_out;
Delay3No1_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_4_cast <= Delay3No1_out;
   MUX_Add11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No66_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg108_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay3No1_out_to_MUX_Add11_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add11_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add4_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add4_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add4_impl_out,
                 X => Delay1No36_out_to_Add4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add4_impl_parent_implementedSystem_port_1_cast);

SharedReg55_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg55_out;
SharedReg4_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg72_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg72_out;
SharedReg101_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
   MUX_Add4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg55_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg72_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Add4_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add4_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add4_impl_0_out,
                 Y => Delay1No36_out);

SharedReg96_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg20_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg78_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg140_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg140_out;
   MUX_Add4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg78_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg140_out_to_MUX_Add4_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add4_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add4_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add6_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add6_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add6_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add6_impl_out,
                 X => Delay1No38_out_to_Add6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add6_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg5_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg94_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg78_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg78_out;
   MUX_Add6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg78_out_to_MUX_Add6_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add6_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_impl_0_out,
                 Y => Delay1No38_out);

SharedReg72_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg21_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg57_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg85_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg85_out;
   MUX_Add6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg85_out_to_MUX_Add6_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add6_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add6_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add15_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add15_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add15_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add15_impl_out,
                 X => Delay1No40_out_to_Add15_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add15_impl_parent_implementedSystem_port_1_cast);

SharedReg103_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast <= SharedReg103_out;
SharedReg12_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg67_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg88_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_4_cast <= SharedReg88_out;
   MUX_Add15_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg103_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg67_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg88_out_to_MUX_Add15_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add15_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_impl_0_out,
                 Y => Delay1No40_out);

SharedReg51_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast <= SharedReg51_out;
SharedReg28_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg93_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_3_cast <= SharedReg93_out;
SharedReg108_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_4_cast <= SharedReg108_out;
   MUX_Add15_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg51_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg93_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg108_out_to_MUX_Add15_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add15_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add15_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add7_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add7_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add7_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add7_impl_out,
                 X => Delay1No42_out_to_Add7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add7_impl_parent_implementedSystem_port_1_cast);

SharedReg120_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg120_out;
SharedReg78_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg78_out;
SharedReg95_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg51_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg51_out;
   MUX_Add7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg120_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg51_out_to_MUX_Add7_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add7_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_0_out,
                 Y => Delay1No42_out);

SharedReg67_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg67_out;
SharedReg93_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg93_out;
SharedReg102_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg102_out;
SharedReg55_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg55_out;
   MUX_Add7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg67_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg102_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg55_out_to_MUX_Add7_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add7_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add7_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add16_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add16_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add16_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add16_impl_out,
                 X => Delay1No44_out_to_Add16_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add16_impl_parent_implementedSystem_port_1_cast);

SharedReg104_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg60_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast <= SharedReg60_out;
SharedReg85_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_3_cast <= SharedReg85_out;
SharedReg93_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_4_cast <= SharedReg93_out;
   MUX_Add16_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg60_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg85_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg93_out_to_MUX_Add16_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_impl_0_out,
                 Y => Delay1No44_out);

SharedReg52_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast <= SharedReg52_out;
SharedReg61_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg101_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_3_cast <= SharedReg101_out;
SharedReg110_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_4_cast <= SharedReg110_out;
   MUX_Add16_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg52_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg101_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Add16_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add16_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add16_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add9_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add9_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add9_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_impl_out,
                 X => Delay1No46_out_to_Add9_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add9_impl_parent_implementedSystem_port_1_cast);

SharedReg73_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg110_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast <= SharedReg110_out;
SharedReg103_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg52_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_4_cast <= SharedReg52_out;
   MUX_Add9_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg52_out_to_MUX_Add9_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add9_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_0_out,
                 Y => Delay1No46_out);

SharedReg78_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg113_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast <= SharedReg113_out;
SharedReg125_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg56_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_4_cast <= SharedReg56_out;
   MUX_Add9_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg113_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg125_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_Add9_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add9_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add18_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add18_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add18_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_impl_out,
                 X => Delay1No48_out_to_Add18_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add18_impl_parent_implementedSystem_port_1_cast);

SharedReg50_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast <= SharedReg50_out;
SharedReg103_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast <= SharedReg103_out;
SharedReg104_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_3_cast <= SharedReg104_out;
SharedReg113_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_4_cast <= SharedReg113_out;
   MUX_Add18_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg50_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg103_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg104_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg113_out_to_MUX_Add18_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add18_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_0_out,
                 Y => Delay1No48_out);

SharedReg53_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg104_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast <= SharedReg104_out;
SharedReg126_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_3_cast <= SharedReg126_out;
SharedReg69_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_4_cast <= SharedReg69_out;
   MUX_Add18_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg126_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg69_out_to_MUX_Add18_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add18_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add111_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add111_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add111_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_impl_out,
                 X => Delay1No50_out_to_Add111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add111_impl_parent_implementedSystem_port_1_cast);

SharedReg93_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast <= SharedReg93_out;
SharedReg85_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg85_out;
Delay2No4_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_3_cast <= Delay2No4_out;
SharedReg58_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_4_cast <= SharedReg58_out;
   MUX_Add111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg93_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg85_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No4_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg58_out_to_MUX_Add111_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add111_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_impl_0_out,
                 Y => Delay1No50_out);

SharedReg85_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg85_out;
SharedReg88_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast <= SharedReg88_out;
Delay2No13_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_3_cast <= Delay2No13_out;
SharedReg59_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_4_cast <= SharedReg59_out;
   MUX_Add111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg85_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg88_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No13_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg59_out_to_MUX_Add111_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add111_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add22_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add22_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add22_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add22_impl_out,
                 X => Delay1No52_out_to_Add22_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add22_impl_parent_implementedSystem_port_1_cast);

SharedReg56_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg62_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg11_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg118_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_4_cast <= SharedReg118_out;
   MUX_Add22_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg11_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg118_out_to_MUX_Add22_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add22_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_impl_0_out,
                 Y => Delay1No52_out);

SharedReg58_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast <= SharedReg58_out;
SharedReg94_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast <= SharedReg94_out;
SharedReg27_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg120_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_4_cast <= SharedReg120_out;
   MUX_Add22_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg58_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg27_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg120_out_to_MUX_Add22_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add22_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add22_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add112_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add112_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add112_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add112_impl_out,
                 X => Delay1No54_out_to_Add112_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add112_impl_parent_implementedSystem_port_1_cast);

SharedReg60_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg101_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast <= SharedReg101_out;
SharedReg64_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_3_cast <= SharedReg64_out;
SharedReg60_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
   MUX_Add112_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg64_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Add112_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add112_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add112_impl_0_out,
                 Y => Delay1No54_out);

SharedReg61_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg108_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast <= SharedReg108_out;
SharedReg65_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_3_cast <= SharedReg65_out;
SharedReg61_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_4_cast <= SharedReg61_out;
   MUX_Add112_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg65_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg61_out_to_MUX_Add112_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add112_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add112_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add121_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add121_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add121_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add121_impl_out,
                 X => Delay1No56_out_to_Add121_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add121_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg95_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg75_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_3_cast <= SharedReg75_out;
SharedReg47_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_4_cast <= SharedReg47_out;
   MUX_Add121_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg75_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg47_out_to_MUX_Add121_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add121_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_impl_0_out,
                 Y => Delay1No56_out);

SharedReg101_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg102_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_2_cast <= SharedReg102_out;
SharedReg76_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_3_cast <= SharedReg76_out;
SharedReg62_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
   MUX_Add121_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg102_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg76_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Add121_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add121_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add121_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add33_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add33_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add33_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add33_impl_out,
                 X => Delay1No58_out_to_Add33_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add33_impl_parent_implementedSystem_port_1_cast);

SharedReg62_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_1_cast <= SharedReg62_out;
SharedReg118_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
SharedReg82_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_3_cast <= SharedReg82_out;
SharedReg63_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_4_cast <= SharedReg63_out;
   MUX_Add33_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg62_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg82_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg63_out_to_MUX_Add33_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add33_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_impl_0_out,
                 Y => Delay1No58_out);

SharedReg94_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg120_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_2_cast <= SharedReg120_out;
SharedReg83_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_3_cast <= SharedReg83_out;
SharedReg64_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_4_cast <= SharedReg64_out;
   MUX_Add33_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg120_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg83_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg64_out_to_MUX_Add33_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add33_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add33_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add34_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add34_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add34_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add34_impl_out,
                 X => Delay1No60_out_to_Add34_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add34_impl_parent_implementedSystem_port_1_cast);

SharedReg108_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_1_cast <= SharedReg108_out;
SharedReg6_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg71_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_3_cast <= SharedReg71_out;
SharedReg65_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_4_cast <= SharedReg65_out;
   MUX_Add34_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg108_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg71_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg65_out_to_MUX_Add34_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add34_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add34_impl_0_out,
                 Y => Delay1No60_out);

SharedReg110_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_1_cast <= SharedReg110_out;
SharedReg22_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
Delay2No43_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_3_cast <= Delay2No43_out;
SharedReg66_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_4_cast <= SharedReg66_out;
   MUX_Add34_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg110_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No43_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg66_out_to_MUX_Add34_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add34_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add34_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add124_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add124_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add124_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add124_impl_out,
                 X => Delay1No62_out_to_Add124_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add124_impl_parent_implementedSystem_port_1_cast);

SharedReg95_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_1_cast <= SharedReg95_out;
SharedReg7_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg90_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg76_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_4_cast <= SharedReg76_out;
   MUX_Add124_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg95_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg90_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg76_out_to_MUX_Add124_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add124_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add124_impl_0_out,
                 Y => Delay1No62_out);

SharedReg102_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_1_cast <= SharedReg102_out;
SharedReg23_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg91_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_3_cast <= SharedReg91_out;
SharedReg77_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_4_cast <= SharedReg77_out;
   MUX_Add124_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg102_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg91_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg77_out_to_MUX_Add124_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add124_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add124_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add37_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add37_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add37_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add37_impl_out,
                 X => Delay1No64_out_to_Add37_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add37_impl_parent_implementedSystem_port_1_cast);

SharedReg68_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_1_cast <= SharedReg68_out;
SharedReg8_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg98_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg81_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_4_cast <= SharedReg81_out;
   MUX_Add37_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg68_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg98_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg81_out_to_MUX_Add37_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add37_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add37_impl_0_out,
                 Y => Delay1No64_out);

Delay2No60_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_1_cast <= Delay2No60_out;
SharedReg24_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg99_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg82_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_4_cast <= SharedReg82_out;
   MUX_Add37_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No60_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg99_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg82_out_to_MUX_Add37_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add37_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add37_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add127_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add127_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add127_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add127_impl_out,
                 X => Delay1No66_out_to_Add127_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add127_impl_parent_implementedSystem_port_1_cast);

SharedReg63_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_1_cast <= SharedReg63_out;
SharedReg9_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_2_cast <= SharedReg9_out;
SharedReg105_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_3_cast <= SharedReg105_out;
Delay2No56_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_4_cast <= Delay2No56_out;
   MUX_Add127_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg63_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg9_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg105_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No56_out_to_MUX_Add127_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add127_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_impl_0_out,
                 Y => Delay1No66_out);

SharedReg64_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_1_cast <= SharedReg64_out;
SharedReg25_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_2_cast <= SharedReg25_out;
Delay2No48_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_3_cast <= Delay2No48_out;
SharedReg84_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_4_cast <= SharedReg84_out;
   MUX_Add127_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg64_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg25_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No48_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg84_out_to_MUX_Add127_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add127_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add127_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add129_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add129_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add129_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add129_impl_out,
                 X => Delay1No68_out_to_Add129_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add129_impl_parent_implementedSystem_port_1_cast);

SharedReg65_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg13_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg107_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_3_cast <= SharedReg107_out;
SharedReg97_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_4_cast <= SharedReg97_out;
   MUX_Add129_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg107_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg97_out_to_MUX_Add129_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add129_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_impl_0_out,
                 Y => Delay1No68_out);

SharedReg66_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_1_cast <= SharedReg66_out;
SharedReg29_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg109_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_3_cast <= SharedReg109_out;
SharedReg98_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_4_cast <= SharedReg98_out;
   MUX_Add129_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg66_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg109_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg98_out_to_MUX_Add129_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add129_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add129_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add40_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add40_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add40_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_impl_out,
                 X => Delay1No70_out_to_Add40_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add40_impl_parent_implementedSystem_port_1_cast);

SharedReg81_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_1_cast <= SharedReg81_out;
SharedReg14_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_2_cast <= SharedReg14_out;
Delay3No3_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_3_cast <= Delay3No3_out;
SharedReg105_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_4_cast <= SharedReg105_out;
   MUX_Add40_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg81_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg14_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No3_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg105_out_to_MUX_Add40_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add40_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_impl_0_out,
                 Y => Delay1No70_out);

SharedReg82_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_1_cast <= SharedReg82_out;
SharedReg30_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_2_cast <= SharedReg30_out;
Delay2No52_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_3_cast <= Delay2No52_out;
SharedReg106_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_4_cast <= SharedReg106_out;
   MUX_Add40_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg82_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg30_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No52_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg106_out_to_MUX_Add40_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add40_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add130_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add130_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add130_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add130_impl_out,
                 X => Delay1No72_out_to_Add130_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add130_impl_parent_implementedSystem_port_1_cast);

SharedReg87_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_1_cast <= SharedReg87_out;
SharedReg15_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg115_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg109_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_4_cast <= SharedReg109_out;
   MUX_Add130_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg87_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg115_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg109_out_to_MUX_Add130_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add130_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_impl_0_out,
                 Y => Delay1No72_out);

SharedReg89_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg31_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg116_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_3_cast <= SharedReg116_out;
SharedReg111_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_4_cast <= SharedReg111_out;
   MUX_Add130_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg116_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg111_out_to_MUX_Add130_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add130_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add130_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add42_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add42_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add42_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add42_impl_out,
                 X => Delay1No74_out_to_Add42_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add42_impl_parent_implementedSystem_port_1_cast);

SharedReg76_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_1_cast <= SharedReg76_out;
SharedReg72_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
Delay2No54_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_3_cast <= Delay2No54_out;
SharedReg112_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_4_cast <= SharedReg112_out;
   MUX_Add42_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg76_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No54_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg112_out_to_MUX_Add42_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add42_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add42_impl_0_out,
                 Y => Delay1No74_out);

SharedReg77_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_1_cast <= SharedReg77_out;
SharedReg114_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_2_cast <= SharedReg114_out;
SharedReg119_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_3_cast <= SharedReg119_out;
SharedReg115_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_4_cast <= SharedReg115_out;
   MUX_Add42_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg77_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg119_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg115_out_to_MUX_Add42_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add42_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add42_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add1_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add1_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add1_impl_out,
                 X => Delay1No76_out_to_Add1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add1_impl_parent_implementedSystem_port_1_cast);

SharedReg97_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg55_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg55_out;
SharedReg128_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg128_out;
SharedReg89_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg89_out;
   MUX_Add1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg128_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg89_out_to_MUX_Add1_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add1_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add1_impl_0_out,
                 Y => Delay1No76_out);

SharedReg98_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg98_out;
SharedReg125_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg125_out;
SharedReg129_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg129_out;
SharedReg90_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg90_out;
   MUX_Add1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg125_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg129_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg90_out_to_MUX_Add1_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add1_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add1_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product4_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product4_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_impl_out,
                 X => Delay1No78_out_to_Product4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product4_impl_parent_implementedSystem_port_1_cast);

SharedReg164_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg179_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg179_out;
SharedReg162_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg162_out;
Delay7No1_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_4_cast <= Delay7No1_out;
   MUX_Product4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg179_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg162_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay7No1_out_to_MUX_Product4_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product4_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_0_out,
                 Y => Delay1No78_out);

SharedReg33_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg33_out;
SharedReg53_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg53_out;
SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg153_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg153_out;
   MUX_Product4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg33_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg53_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg153_out_to_MUX_Product4_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product4_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product11_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product11_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product11_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_impl_out,
                 X => Delay1No80_out_to_Product11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product11_impl_parent_implementedSystem_port_1_cast);

Delay8No2_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast <= Delay8No2_out;
SharedReg49_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg49_out;
SharedReg162_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_3_cast <= SharedReg162_out;
Delay7No2_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_4_cast <= Delay7No2_out;
   MUX_Product11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay8No2_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg49_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg162_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay7No2_out_to_MUX_Product11_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_impl_0_out,
                 Y => Delay1No80_out);

SharedReg34_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast <= SharedReg34_out;
SharedReg179_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg179_out;
SharedReg34_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_3_cast <= SharedReg34_out;
Delay2No76_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_4_cast <= Delay2No76_out;
   MUX_Product11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg34_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg179_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg34_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No76_out_to_MUX_Product11_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product11_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product21_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product21_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product21_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_impl_out,
                 X => Delay1No82_out_to_Product21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product21_impl_parent_implementedSystem_port_1_cast);

SharedReg188_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast <= SharedReg188_out;
SharedReg197_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast <= SharedReg197_out;
SharedReg163_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_3_cast <= SharedReg163_out;
Delay7No3_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_4_cast <= Delay7No3_out;
   MUX_Product21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg188_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg197_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg163_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay7No3_out_to_MUX_Product21_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product21_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_0_out,
                 Y => Delay1No82_out);

SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg37_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast <= SharedReg37_out;
SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg158_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_4_cast <= SharedReg158_out;
   MUX_Product21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg37_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg158_out_to_MUX_Product21_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product21_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product31_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product31_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product31_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_impl_out,
                 X => Delay1No84_out_to_Product31_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product31_impl_parent_implementedSystem_port_1_cast);

SharedReg189_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast <= SharedReg189_out;
SharedReg32_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast <= SharedReg32_out;
SharedReg34_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_3_cast <= SharedReg34_out;
SharedReg171_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_4_cast <= SharedReg171_out;
   MUX_Product31_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg189_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg34_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg171_out_to_MUX_Product31_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product31_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_impl_0_out,
                 Y => Delay1No84_out);

SharedReg38_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg197_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast <= SharedReg197_out;
SharedReg163_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_3_cast <= SharedReg163_out;
SharedReg155_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_4_cast <= SharedReg155_out;
   MUX_Product31_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg197_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg163_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg155_out_to_MUX_Product31_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product31_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Subtract2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_impl_out,
                 X => Delay1No86_out_to_Subtract2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Subtract2_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg79_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg79_out;
SharedReg63_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg63_out;
SharedReg75_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg75_out;
   MUX_Subtract2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg79_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg63_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg75_out_to_MUX_Subtract2_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract2_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_0_out,
                 Y => Delay1No86_out);

SharedReg83_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg83_out;
SharedReg82_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg66_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg66_out;
SharedReg79_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg79_out;
   MUX_Subtract2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg83_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg66_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg79_out_to_MUX_Subtract2_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract2_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product5_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product5_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_impl_out,
                 X => Delay1No88_out_to_Product5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product5_impl_parent_implementedSystem_port_1_cast);

SharedReg164_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg164_out;
SharedReg178_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg178_out;
SharedReg152_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg152_out;
SharedReg32_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg32_out;
   MUX_Product5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg164_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg178_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg152_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product5_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product5_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_impl_0_out,
                 Y => Delay1No88_out);

SharedReg34_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg34_out;
SharedReg49_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg49_out;
SharedReg169_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg169_out;
SharedReg165_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg165_out;
   MUX_Product5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg34_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg49_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg169_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg165_out_to_MUX_Product5_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product5_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Subtract3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract3_impl_out,
                 X => Delay1No90_out_to_Subtract3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Subtract3_impl_parent_implementedSystem_port_1_cast);

SharedReg70_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg74_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg74_out;
SharedReg79_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg79_out;
Delay2No39_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_4_cast <= Delay2No39_out;
   MUX_Subtract3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg74_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg79_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No39_out_to_MUX_Subtract3_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_impl_0_out,
                 Y => Delay1No90_out);

SharedReg71_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg71_out;
SharedReg77_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg77_out;
SharedReg70_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg70_out;
SharedReg74_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg74_out;
   MUX_Subtract3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg71_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg77_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg70_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg74_out_to_MUX_Subtract3_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract3_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract3_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product6_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product6_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product6_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_impl_out,
                 X => Delay1No92_out_to_Product6_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product6_impl_parent_implementedSystem_port_1_cast);

SharedReg196_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast <= SharedReg196_out;
SharedReg182_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast <= SharedReg182_out;
SharedReg166_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_3_cast <= SharedReg166_out;
SharedReg158_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_4_cast <= SharedReg158_out;
   MUX_Product6_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg196_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg166_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg158_out_to_MUX_Product6_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product6_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_impl_0_out,
                 Y => Delay1No92_out);

SharedReg36_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg38_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg142_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg171_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_4_cast <= SharedReg171_out;
   MUX_Product6_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg171_out_to_MUX_Product6_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product6_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product13_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product13_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product13_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product13_impl_out,
                 X => Delay1No94_out_to_Product13_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product13_impl_parent_implementedSystem_port_1_cast);

SharedReg216_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast <= SharedReg216_out;
SharedReg182_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast <= SharedReg182_out;
SharedReg166_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_3_cast <= SharedReg166_out;
SharedReg172_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_4_cast <= SharedReg172_out;
   MUX_Product13_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg216_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg182_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg166_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg172_out_to_MUX_Product13_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product13_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_0_out,
                 Y => Delay1No94_out);

SharedReg41_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg39_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg145_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_3_cast <= SharedReg145_out;
SharedReg157_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_4_cast <= SharedReg157_out;
   MUX_Product13_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg145_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg157_out_to_MUX_Product13_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product13_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product13_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product23_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product23_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product23_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_impl_out,
                 X => Delay1No96_out_to_Product23_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product23_impl_parent_implementedSystem_port_1_cast);

SharedReg216_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast <= SharedReg216_out;
SharedReg183_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast <= SharedReg183_out;
SharedReg167_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_3_cast <= SharedReg167_out;
SharedReg172_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_4_cast <= SharedReg172_out;
   MUX_Product23_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg216_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg183_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg167_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg172_out_to_MUX_Product23_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product23_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_0_out,
                 Y => Delay1No96_out);

SharedReg42_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg38_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg142_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg159_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_4_cast <= SharedReg159_out;
   MUX_Product23_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product23_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product23_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product33_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product33_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product33_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_impl_out,
                 X => Delay1No98_out_to_Product33_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product33_impl_parent_implementedSystem_port_1_cast);

SharedReg217_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast <= SharedReg217_out;
SharedReg39_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg145_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_3_cast <= SharedReg145_out;
SharedReg173_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_4_cast <= SharedReg173_out;
   MUX_Product33_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg217_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg145_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg173_out_to_MUX_Product33_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product33_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_0_out,
                 Y => Delay1No98_out);

SharedReg41_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast <= SharedReg41_out;
SharedReg183_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast <= SharedReg183_out;
SharedReg167_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_3_cast <= SharedReg167_out;
SharedReg157_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_4_cast <= SharedReg157_out;
   MUX_Product33_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg41_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg183_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg167_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg157_out_to_MUX_Product33_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product33_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Subtract4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_impl_out,
                 X => Delay1No100_out_to_Subtract4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Subtract4_impl_parent_implementedSystem_port_1_cast);

SharedReg84_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg83_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg83_out;
SharedReg74_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg80_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg80_out;
   MUX_Subtract4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg83_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg74_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg80_out_to_MUX_Subtract4_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract4_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_0_out,
                 Y => Delay1No100_out);

SharedReg90_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg84_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg84_out;
SharedReg77_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg77_out;
SharedReg83_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg83_out;
   MUX_Subtract4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg84_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg77_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg83_out_to_MUX_Subtract4_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract4_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product7_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product7_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product7_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product7_impl_out,
                 X => Delay1No102_out_to_Product7_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product7_impl_parent_implementedSystem_port_1_cast);

SharedReg200_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast <= SharedReg200_out;
SharedReg184_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast <= SharedReg184_out;
SharedReg168_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_3_cast <= SharedReg168_out;
SharedReg159_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_4_cast <= SharedReg159_out;
   MUX_Product7_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg200_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg184_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg168_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg159_out_to_MUX_Product7_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product7_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product7_impl_0_out,
                 Y => Delay1No102_out);

SharedReg154_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast <= SharedReg154_out;
SharedReg40_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg151_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg173_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_4_cast <= SharedReg173_out;
   MUX_Product7_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg154_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg151_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg173_out_to_MUX_Product7_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product7_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product7_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product8_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product8_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product8_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product8_impl_out,
                 X => Delay1No104_out_to_Product8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product8_impl_parent_implementedSystem_port_1_cast);

SharedReg212_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg212_out;
SharedReg184_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg184_out;
SharedReg170_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg170_out;
SharedReg176_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg176_out;
   MUX_Product8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg212_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg184_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg170_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg176_out_to_MUX_Product8_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product8_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product8_impl_0_out,
                 Y => Delay1No104_out);

SharedReg124_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg41_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg154_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg154_out;
SharedReg160_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg160_out;
   MUX_Product8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg154_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg160_out_to_MUX_Product8_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product8_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product8_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product10_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product10_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product10_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_impl_out,
                 X => Delay1No106_out_to_Product10_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product10_impl_parent_implementedSystem_port_1_cast);

SharedReg212_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast <= SharedReg212_out;
SharedReg185_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast <= SharedReg185_out;
SharedReg206_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_3_cast <= SharedReg206_out;
SharedReg176_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_4_cast <= SharedReg176_out;
   MUX_Product10_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg212_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg185_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg206_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg176_out_to_MUX_Product10_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product10_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_0_out,
                 Y => Delay1No106_out);

SharedReg131_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg40_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast <= SharedReg40_out;
SharedReg158_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_3_cast <= SharedReg158_out;
SharedReg161_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_4_cast <= SharedReg161_out;
   MUX_Product10_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg40_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg158_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg161_out_to_MUX_Product10_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product10_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product17_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product17_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product17_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product17_impl_out,
                 X => Delay1No108_out_to_Product17_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product17_impl_parent_implementedSystem_port_1_cast);

SharedReg213_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_1_cast <= SharedReg213_out;
SharedReg41_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg206_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_3_cast <= SharedReg206_out;
SharedReg177_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_4_cast <= SharedReg177_out;
   MUX_Product17_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg206_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg177_out_to_MUX_Product17_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product17_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_impl_0_out,
                 Y => Delay1No108_out);

SharedReg124_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_1_cast <= SharedReg124_out;
SharedReg185_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_2_cast <= SharedReg185_out;
SharedReg159_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_3_cast <= SharedReg159_out;
SharedReg160_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_4_cast <= SharedReg160_out;
   MUX_Product17_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg124_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg185_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg159_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg160_out_to_MUX_Product17_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product17_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product17_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product27_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product27_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product27_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product27_impl_out,
                 X => Delay1No110_out_to_Product27_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product27_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
Delay21No14_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_2_cast <= Delay21No14_out;
SharedReg207_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_3_cast <= SharedReg207_out;
SharedReg161_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_4_cast <= SharedReg161_out;
   MUX_Product27_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay21No14_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg207_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg161_out_to_MUX_Product27_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_impl_0_out,
                 Y => Delay1No110_out);

SharedReg213_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_1_cast <= SharedReg213_out;
Delay2No24_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_2_cast <= Delay2No24_out;
SharedReg158_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_3_cast <= SharedReg158_out;
SharedReg177_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_4_cast <= SharedReg177_out;
   MUX_Product27_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay2No24_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg158_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg177_out_to_MUX_Product27_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product27_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product27_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product37_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product37_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product37_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_impl_out,
                 X => Delay1No112_out_to_Product37_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product37_impl_parent_implementedSystem_port_1_cast);

SharedReg214_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast <= SharedReg214_out;
SharedReg33_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast <= SharedReg33_out;
SharedReg159_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_3_cast <= SharedReg159_out;
Delay7No14_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_4_cast <= Delay7No14_out;
   MUX_Product37_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg214_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg33_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg159_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay7No14_out_to_MUX_Product37_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product37_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_impl_0_out,
                 Y => Delay1No112_out);

SharedReg39_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
Delay21No15_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast <= Delay21No15_out;
SharedReg207_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_3_cast <= SharedReg207_out;
Delay2No27_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_4_cast <= Delay2No27_out;
   MUX_Product37_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay21No15_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg207_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No27_out_to_MUX_Product37_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product37_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Subtract8_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Subtract8_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Subtract8_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract8_impl_out,
                 X => Delay1No114_out_to_Subtract8_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Subtract8_impl_parent_implementedSystem_port_1_cast);

SharedReg92_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg92_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_2_cast <= SharedReg92_out;
SharedReg81_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_3_cast <= SharedReg81_out;
SharedReg100_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_4_cast <= SharedReg100_out;
   MUX_Subtract8_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg92_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg81_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg100_out_to_MUX_Subtract8_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract8_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_impl_0_out,
                 Y => Delay1No114_out);

SharedReg99_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_1_cast <= SharedReg99_out;
SharedReg99_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_2_cast <= SharedReg99_out;
SharedReg84_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg107_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_4_cast <= SharedReg107_out;
   MUX_Subtract8_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg99_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg99_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg84_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg107_out_to_MUX_Subtract8_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract8_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract8_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product20_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product20_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product20_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product20_impl_out,
                 X => Delay1No116_out_to_Product20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product20_impl_parent_implementedSystem_port_1_cast);

SharedReg214_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_1_cast <= SharedReg214_out;
SharedReg190_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_2_cast <= SharedReg190_out;
Delay22No1_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_3_cast <= Delay22No1_out;
SharedReg240_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_4_cast <= SharedReg240_out;
   MUX_Product20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg214_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg190_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No1_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg240_out_to_MUX_Product20_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product20_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product20_impl_0_out,
                 Y => Delay1No116_out);

SharedReg40_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg42_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg54_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_3_cast <= SharedReg54_out;
SharedReg41_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_4_cast <= SharedReg41_out;
   MUX_Product20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg54_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg41_out_to_MUX_Product20_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product20_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product20_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Subtract10_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Subtract10_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Subtract10_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract10_impl_out,
                 X => Delay1No118_out_to_Subtract10_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Subtract10_impl_parent_implementedSystem_port_1_cast);

SharedReg100_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_1_cast <= SharedReg100_out;
SharedReg100_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg87_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_3_cast <= SharedReg87_out;
SharedReg87_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_4_cast <= SharedReg87_out;
   MUX_Subtract10_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg100_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg87_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg87_out_to_MUX_Subtract10_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract10_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_impl_0_out,
                 Y => Delay1No118_out);

SharedReg107_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg107_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_2_cast <= SharedReg107_out;
Delay2No44_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_3_cast <= Delay2No44_out;
SharedReg91_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_4_cast <= SharedReg91_out;
   MUX_Subtract10_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg107_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No44_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg91_out_to_MUX_Subtract10_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract10_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract10_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product30_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product30_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product30_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product30_impl_out,
                 X => Delay1No120_out_to_Product30_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product30_impl_parent_implementedSystem_port_1_cast);

SharedReg215_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg190_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_2_cast <= SharedReg190_out;
SharedReg180_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_3_cast <= SharedReg180_out;
SharedReg240_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_4_cast <= SharedReg240_out;
   MUX_Product30_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg190_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg180_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg240_out_to_MUX_Product30_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product30_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product30_impl_0_out,
                 Y => Delay1No120_out);

SharedReg39_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg43_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg61_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_3_cast <= SharedReg61_out;
SharedReg42_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_4_cast <= SharedReg42_out;
   MUX_Product30_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg61_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg42_out_to_MUX_Product30_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product30_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product30_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product111_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product111_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product111_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_impl_out,
                 X => Delay1No122_out_to_Product111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product111_impl_parent_implementedSystem_port_1_cast);

SharedReg40_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast <= SharedReg40_out;
SharedReg191_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg191_out;
SharedReg180_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_3_cast <= SharedReg180_out;
SharedReg241_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_4_cast <= SharedReg241_out;
   MUX_Product111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg40_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg180_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_Product111_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_0_out,
                 Y => Delay1No122_out);

SharedReg215_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg42_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast <= SharedReg42_out;
SharedReg62_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg41_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_4_cast <= SharedReg41_out;
   MUX_Product111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg42_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg62_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg41_out_to_MUX_Product111_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product111_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product210_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product210_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product210_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_impl_out,
                 X => Delay1No124_out_to_Product210_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product210_impl_parent_implementedSystem_port_1_cast);

SharedReg42_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg43_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast <= SharedReg43_out;
SharedReg181_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_3_cast <= SharedReg181_out;
SharedReg42_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_4_cast <= SharedReg42_out;
   MUX_Product210_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg43_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg181_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg42_out_to_MUX_Product210_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_0_out,
                 Y => Delay1No124_out);

SharedReg217_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast <= SharedReg217_out;
SharedReg191_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast <= SharedReg191_out;
SharedReg61_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_3_cast <= SharedReg61_out;
SharedReg241_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_4_cast <= SharedReg241_out;
   MUX_Product210_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg217_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg191_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg61_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg241_out_to_MUX_Product210_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product210_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product310_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product310_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product310_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_impl_out,
                 X => Delay1No126_out_to_Product310_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product310_impl_parent_implementedSystem_port_1_cast);

SharedReg220_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast <= SharedReg220_out;
SharedReg192_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast <= SharedReg192_out;
SharedReg62_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_3_cast <= SharedReg62_out;
SharedReg228_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_4_cast <= SharedReg228_out;
   MUX_Product310_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg220_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg192_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg62_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg228_out_to_MUX_Product310_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_0_out,
                 Y => Delay1No126_out);

SharedReg43_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast <= SharedReg43_out;
SharedReg131_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast <= SharedReg131_out;
SharedReg181_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_3_cast <= SharedReg181_out;
SharedReg36_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
   MUX_Product310_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg43_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg131_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg181_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product310_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product310_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Subtract11_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract11_impl_out,
                 X => Delay1No128_out_to_Subtract11_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Subtract11_impl_parent_implementedSystem_port_1_cast);

SharedReg75_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast <= SharedReg75_out;
SharedReg87_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast <= SharedReg87_out;
SharedReg89_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_3_cast <= SharedReg89_out;
SharedReg92_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_4_cast <= SharedReg92_out;
   MUX_Subtract11_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg75_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg87_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg89_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Subtract11_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract11_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_impl_0_out,
                 Y => Delay1No128_out);

SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast <= SharedReg91_out;
SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast <= SharedReg91_out;
SharedReg92_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_3_cast <= SharedReg92_out;
SharedReg99_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_4_cast <= SharedReg99_out;
   MUX_Subtract11_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg91_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg92_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg99_out_to_MUX_Subtract11_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract11_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract11_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Add53_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Add53_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Add53_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add53_impl_out,
                 X => Delay1No130_out_to_Add53_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Add53_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg75_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_2_cast <= SharedReg75_out;
SharedReg133_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_3_cast <= SharedReg133_out;
SharedReg117_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_4_cast <= SharedReg117_out;
   MUX_Add53_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg75_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg133_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg117_out_to_MUX_Add53_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add53_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add53_impl_0_out,
                 Y => Delay1No130_out);

SharedReg106_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg76_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_2_cast <= SharedReg76_out;
SharedReg134_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_3_cast <= SharedReg134_out;
SharedReg119_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_4_cast <= SharedReg119_out;
   MUX_Add53_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg134_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg119_out_to_MUX_Add53_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add53_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add53_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Add54_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Add54_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Add54_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add54_impl_out,
                 X => Delay1No132_out_to_Add54_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Add54_impl_parent_implementedSystem_port_1_cast);

SharedReg111_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_1_cast <= SharedReg111_out;
SharedReg80_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_2_cast <= SharedReg80_out;
SharedReg137_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_3_cast <= SharedReg137_out;
SharedReg123_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_4_cast <= SharedReg123_out;
   MUX_Add54_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg111_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg80_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg137_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg123_out_to_MUX_Add54_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add54_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_impl_0_out,
                 Y => Delay1No132_out);

SharedReg112_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_1_cast <= SharedReg112_out;
SharedReg81_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_2_cast <= SharedReg81_out;
SharedReg138_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_3_cast <= SharedReg138_out;
SharedReg127_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_4_cast <= SharedReg127_out;
   MUX_Add54_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg112_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg81_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg138_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg127_out_to_MUX_Add54_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Add54_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add54_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product42_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product42_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product42_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product42_impl_out,
                 X => Delay1No134_out_to_Product42_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product42_impl_parent_implementedSystem_port_1_cast);

SharedReg220_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_1_cast <= SharedReg220_out;
SharedReg192_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_2_cast <= SharedReg192_out;
SharedReg186_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_3_cast <= SharedReg186_out;
SharedReg228_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_4_cast <= SharedReg228_out;
   MUX_Product42_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg220_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg192_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg186_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg228_out_to_MUX_Product42_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product42_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_impl_0_out,
                 Y => Delay1No134_out);

SharedReg44_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg140_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_2_cast <= SharedReg140_out;
SharedReg36_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg38_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_4_cast <= SharedReg38_out;
   MUX_Product42_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg140_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg38_out_to_MUX_Product42_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product42_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product42_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product114_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product114_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product114_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product114_impl_out,
                 X => Delay1No136_out_to_Product114_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product114_impl_parent_implementedSystem_port_1_cast);

SharedReg221_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg193_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_2_cast <= SharedReg193_out;
SharedReg186_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_3_cast <= SharedReg186_out;
SharedReg229_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_4_cast <= SharedReg229_out;
   MUX_Product114_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg193_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg186_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg229_out_to_MUX_Product114_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_impl_0_out,
                 Y => Delay1No136_out);

SharedReg43_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_1_cast <= SharedReg43_out;
SharedReg131_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_2_cast <= SharedReg131_out;
SharedReg38_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg36_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_4_cast <= SharedReg36_out;
   MUX_Product114_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg43_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg131_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg36_out_to_MUX_Product114_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product114_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product114_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product213_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product213_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product213_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_impl_out,
                 X => Delay1No138_out_to_Product213_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product213_impl_parent_implementedSystem_port_1_cast);

SharedReg44_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg140_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_2_cast <= SharedReg140_out;
SharedReg187_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_3_cast <= SharedReg187_out;
SharedReg38_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_4_cast <= SharedReg38_out;
   MUX_Product213_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg140_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg187_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg38_out_to_MUX_Product213_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product213_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_impl_0_out,
                 Y => Delay1No138_out);

SharedReg221_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg193_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_2_cast <= SharedReg193_out;
SharedReg36_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg229_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_4_cast <= SharedReg229_out;
   MUX_Product213_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg193_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg229_out_to_MUX_Product213_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product213_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product313_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product313_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product313_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product313_impl_out,
                 X => Delay1No140_out_to_Product313_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product313_impl_parent_implementedSystem_port_1_cast);

SharedReg222_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_1_cast <= SharedReg222_out;
SharedReg194_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_2_cast <= SharedReg194_out;
SharedReg38_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg234_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_4_cast <= SharedReg234_out;
   MUX_Product313_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg222_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg194_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg234_out_to_MUX_Product313_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product313_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_impl_0_out,
                 Y => Delay1No140_out);

SharedReg46_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg142_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_2_cast <= SharedReg142_out;
SharedReg187_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_3_cast <= SharedReg187_out;
SharedReg39_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_4_cast <= SharedReg39_out;
   MUX_Product313_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg142_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg187_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg39_out_to_MUX_Product313_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product313_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product313_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Subtract14_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Subtract14_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Subtract14_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract14_impl_out,
                 X => Delay1No142_out_to_Subtract14_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Subtract14_impl_parent_implementedSystem_port_1_cast);

SharedReg109_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_1_cast <= SharedReg109_out;
SharedReg119_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_2_cast <= SharedReg119_out;
SharedReg97_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_3_cast <= SharedReg97_out;
SharedReg116_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_4_cast <= SharedReg116_out;
   MUX_Subtract14_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg109_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg119_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg97_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg116_out_to_MUX_Subtract14_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract14_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract14_impl_0_out,
                 Y => Delay1No142_out);

SharedReg115_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_1_cast <= SharedReg115_out;
SharedReg123_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_2_cast <= SharedReg123_out;
SharedReg100_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_3_cast <= SharedReg100_out;
SharedReg121_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_4_cast <= SharedReg121_out;
   MUX_Subtract14_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg115_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg100_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg121_out_to_MUX_Subtract14_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract14_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract14_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Add57_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Add57_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Add57_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add57_impl_out,
                 X => Delay1No144_out_to_Add57_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Add57_impl_parent_implementedSystem_port_1_cast);

SharedReg89_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_1_cast <= SharedReg89_out;
SharedReg117_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_2_cast <= SharedReg117_out;
SharedReg130_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_3_cast <= SharedReg130_out;
   MUX_Add57_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg89_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg117_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg130_out_to_MUX_Add57_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Add57_impl_0_LUT_out,
                 oMux => MUX_Add57_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add57_impl_0_out,
                 Y => Delay1No144_out);

SharedReg90_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_1_cast <= SharedReg90_out;
SharedReg119_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_2_cast <= SharedReg119_out;
SharedReg132_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_3_cast <= SharedReg132_out;
   MUX_Add57_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg90_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg119_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg132_out_to_MUX_Add57_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Add57_impl_1_LUT_out,
                 oMux => MUX_Add57_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add57_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Add58_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Add58_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Add58_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add58_impl_out,
                 X => Delay1No146_out_to_Add58_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Add58_impl_parent_implementedSystem_port_1_cast);

SharedReg97_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_1_cast <= SharedReg97_out;
SharedReg123_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_2_cast <= SharedReg123_out;
Delay2No67_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_3_cast <= Delay2No67_out;
   MUX_Add58_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg97_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg123_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No67_out_to_MUX_Add58_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Add58_impl_0_LUT_out,
                 oMux => MUX_Add58_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add58_impl_0_out,
                 Y => Delay1No146_out);

SharedReg98_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_1_cast <= SharedReg98_out;
SharedReg127_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_2_cast <= SharedReg127_out;
SharedReg137_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_3_cast <= SharedReg137_out;
   MUX_Add58_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg137_out_to_MUX_Add58_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Add58_impl_1_LUT_out,
                 oMux => MUX_Add58_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add58_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Add59_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Add59_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Add59_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add59_impl_out,
                 X => Delay1No148_out_to_Add59_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Add59_impl_parent_implementedSystem_port_1_cast);

SharedReg105_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg130_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_2_cast <= SharedReg130_out;
SharedReg139_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_3_cast <= SharedReg139_out;
   MUX_Add59_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg139_out_to_MUX_Add59_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Add59_impl_0_LUT_out,
                 oMux => MUX_Add59_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add59_impl_0_out,
                 Y => Delay1No148_out);

SharedReg106_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_1_cast <= SharedReg106_out;
SharedReg132_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_2_cast <= SharedReg132_out;
SharedReg143_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_3_cast <= SharedReg143_out;
   MUX_Add59_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg106_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg132_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg143_out_to_MUX_Add59_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Add59_impl_1_LUT_out,
                 oMux => MUX_Add59_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add59_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product118_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product118_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product118_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product118_impl_out,
                 X => Delay1No150_out_to_Product118_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product118_impl_parent_implementedSystem_port_1_cast);

SharedReg222_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_1_cast <= SharedReg222_out;
SharedReg194_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_2_cast <= SharedReg194_out;
Delay22No6_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_3_cast <= Delay22No6_out;
SharedReg234_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_4_cast <= SharedReg234_out;
   MUX_Product118_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg222_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg194_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No6_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg234_out_to_MUX_Product118_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product118_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product118_impl_0_out,
                 Y => Delay1No150_out);

SharedReg47_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_1_cast <= SharedReg47_out;
SharedReg145_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_2_cast <= SharedReg145_out;
SharedReg33_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_3_cast <= SharedReg33_out;
SharedReg40_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_4_cast <= SharedReg40_out;
   MUX_Product118_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg33_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg40_out_to_MUX_Product118_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product118_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product118_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product217_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product217_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product217_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product217_impl_out,
                 X => Delay1No152_out_to_Product217_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product217_impl_parent_implementedSystem_port_1_cast);

SharedReg223_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_1_cast <= SharedReg223_out;
SharedReg195_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_2_cast <= SharedReg195_out;
SharedReg198_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg235_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_4_cast <= SharedReg235_out;
   MUX_Product217_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg223_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg195_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg198_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg235_out_to_MUX_Product217_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product217_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product217_impl_0_out,
                 Y => Delay1No152_out);

SharedReg46_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg142_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_2_cast <= SharedReg142_out;
SharedReg35_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_3_cast <= SharedReg35_out;
SharedReg39_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_4_cast <= SharedReg39_out;
   MUX_Product217_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg142_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg35_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg39_out_to_MUX_Product217_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product217_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product217_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product317_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product317_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product317_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product317_impl_out,
                 X => Delay1No154_out_to_Product317_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product317_impl_parent_implementedSystem_port_1_cast);

SharedReg47_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_1_cast <= SharedReg47_out;
SharedReg145_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_2_cast <= SharedReg145_out;
SharedReg198_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_3_cast <= SharedReg198_out;
SharedReg40_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_4_cast <= SharedReg40_out;
   MUX_Product317_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg47_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg198_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg40_out_to_MUX_Product317_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product317_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product317_impl_0_out,
                 Y => Delay1No154_out);

SharedReg223_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_1_cast <= SharedReg223_out;
SharedReg195_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_2_cast <= SharedReg195_out;
SharedReg37_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_3_cast <= SharedReg37_out;
SharedReg235_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_4_cast <= SharedReg235_out;
   MUX_Product317_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg223_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg195_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg37_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg235_out_to_MUX_Product317_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product317_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product317_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Subtract19_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Subtract19_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Subtract19_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract19_impl_out,
                 X => Delay1No156_out_to_Subtract19_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Subtract19_impl_parent_implementedSystem_port_1_cast);

SharedReg116_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_1_cast <= SharedReg116_out;
SharedReg127_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_2_cast <= SharedReg127_out;
Delay3No2_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_3_cast <= Delay3No2_out;
SharedReg122_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_4_cast <= SharedReg122_out;
   MUX_Subtract19_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg116_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg127_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No2_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_Subtract19_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract19_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract19_impl_0_out,
                 Y => Delay1No156_out);

SharedReg121_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_1_cast <= SharedReg121_out;
SharedReg130_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_2_cast <= SharedReg130_out;
Delay2No49_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_3_cast <= Delay2No49_out;
SharedReg128_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_4_cast <= SharedReg128_out;
   MUX_Subtract19_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg121_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg130_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No49_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg128_out_to_MUX_Subtract19_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract19_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract19_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product219_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product219_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product219_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product219_impl_out,
                 X => Delay1No158_out_to_Product219_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product219_impl_parent_implementedSystem_port_1_cast);

SharedReg226_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_1_cast <= SharedReg226_out;
SharedReg36_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_2_cast <= SharedReg36_out;
Delay22No9_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_3_cast <= Delay22No9_out;
SharedReg238_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_4_cast <= SharedReg238_out;
   MUX_Product219_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg36_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No9_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg238_out_to_MUX_Product219_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product219_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product219_impl_0_out,
                 Y => Delay1No158_out);

SharedReg148_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_1_cast <= SharedReg148_out;
SharedReg199_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_2_cast <= SharedReg199_out;
SharedReg35_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_3_cast <= SharedReg35_out;
SharedReg148_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_4_cast <= SharedReg148_out;
   MUX_Product219_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg199_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg35_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg148_out_to_MUX_Product219_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product219_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product219_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Subtract20_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_impl_out,
                 X => Delay1No160_out_to_Subtract20_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Subtract20_impl_parent_implementedSystem_port_1_cast);

SharedReg122_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg103_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast <= SharedReg103_out;
SharedReg106_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_3_cast <= SharedReg106_out;
SharedReg129_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_4_cast <= SharedReg129_out;
   MUX_Subtract20_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg103_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg106_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg129_out_to_MUX_Subtract20_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract20_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_impl_0_out,
                 Y => Delay1No160_out);

SharedReg128_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast <= SharedReg128_out;
SharedReg104_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast <= SharedReg104_out;
Delay2No50_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_3_cast <= Delay2No50_out;
SharedReg133_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_4_cast <= SharedReg133_out;
   MUX_Subtract20_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg128_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No50_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg133_out_to_MUX_Subtract20_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract20_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product49_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product49_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product49_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product49_impl_out,
                 X => Delay1No162_out_to_Product49_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product49_impl_parent_implementedSystem_port_1_cast);

SharedReg226_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_1_cast <= SharedReg226_out;
Delay21No31_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_2_cast <= Delay21No31_out;
Delay3No9_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_3_cast <= Delay3No9_out;
SharedReg239_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_4_cast <= SharedReg239_out;
   MUX_Product49_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay21No31_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No9_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg239_out_to_MUX_Product49_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product49_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product49_impl_0_out,
                 Y => Delay1No162_out);

SharedReg149_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg153_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_2_cast <= SharedReg153_out;
Delay22No10_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_3_cast <= Delay22No10_out;
SharedReg147_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_4_cast <= SharedReg147_out;
   MUX_Product49_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No10_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_Product49_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product49_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product49_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product220_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product220_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product220_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product220_impl_out,
                 X => Delay1No164_out_to_Product220_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product220_impl_parent_implementedSystem_port_1_cast);

SharedReg227_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg201_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_2_cast <= SharedReg201_out;
SharedReg202_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_3_cast <= SharedReg202_out;
SharedReg236_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_4_cast <= SharedReg236_out;
   MUX_Product220_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg201_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg202_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg236_out_to_MUX_Product220_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product220_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_impl_0_out,
                 Y => Delay1No164_out);

SharedReg148_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_1_cast <= SharedReg148_out;
SharedReg153_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_2_cast <= SharedReg153_out;
SharedReg160_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_3_cast <= SharedReg160_out;
SharedReg150_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_4_cast <= SharedReg150_out;
   MUX_Product220_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg148_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg153_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg160_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg150_out_to_MUX_Product220_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product220_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Subtract21_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Subtract21_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Subtract21_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract21_impl_out,
                 X => Delay1No166_out_to_Subtract21_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Subtract21_impl_parent_implementedSystem_port_1_cast);

SharedReg129_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_1_cast <= SharedReg129_out;
SharedReg85_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_2_cast <= SharedReg85_out;
Delay2No51_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_3_cast <= Delay2No51_out;
SharedReg134_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_4_cast <= SharedReg134_out;
   MUX_Subtract21_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg129_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg85_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No51_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg134_out_to_MUX_Subtract21_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract21_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_impl_0_out,
                 Y => Delay1No166_out);

SharedReg133_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg88_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_2_cast <= SharedReg88_out;
SharedReg111_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_3_cast <= SharedReg111_out;
SharedReg135_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_4_cast <= SharedReg135_out;
   MUX_Subtract21_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg88_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg111_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg135_out_to_MUX_Subtract21_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract21_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract21_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product122_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product122_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product122_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product122_impl_out,
                 X => Delay1No168_out_to_Product122_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product122_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg174_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_2_cast <= SharedReg174_out;
SharedReg202_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_3_cast <= SharedReg202_out;
SharedReg237_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_4_cast <= SharedReg237_out;
   MUX_Product122_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg202_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg237_out_to_MUX_Product122_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product122_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_impl_0_out,
                 Y => Delay1No168_out);

SharedReg227_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg141_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
SharedReg161_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_3_cast <= SharedReg161_out;
SharedReg149_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_4_cast <= SharedReg149_out;
   MUX_Product122_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg161_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg149_out_to_MUX_Product122_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product122_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product122_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product221_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product221_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product221_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product221_impl_out,
                 X => Delay1No170_out_to_Product221_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product221_impl_parent_implementedSystem_port_1_cast);

SharedReg224_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast <= SharedReg224_out;
SharedReg174_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast <= SharedReg174_out;
SharedReg203_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_3_cast <= SharedReg203_out;
SharedReg242_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_4_cast <= SharedReg242_out;
   MUX_Product221_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg224_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg203_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg242_out_to_MUX_Product221_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product221_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_impl_0_out,
                 Y => Delay1No170_out);

SharedReg150_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast <= SharedReg150_out;
SharedReg124_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast <= SharedReg124_out;
SharedReg160_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_3_cast <= SharedReg160_out;
SharedReg34_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_4_cast <= SharedReg34_out;
   MUX_Product221_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg150_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg160_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg34_out_to_MUX_Product221_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product221_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product221_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product321_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product321_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product321_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product321_impl_out,
                 X => Delay1No172_out_to_Product321_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product321_impl_parent_implementedSystem_port_1_cast);

SharedReg224_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast <= SharedReg224_out;
SharedReg124_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast <= SharedReg124_out;
SharedReg161_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_3_cast <= SharedReg161_out;
SharedReg242_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_4_cast <= SharedReg242_out;
   MUX_Product321_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg224_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg124_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg161_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg242_out_to_MUX_Product321_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product321_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_0_out,
                 Y => Delay1No172_out);

SharedReg151_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg175_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast <= SharedReg175_out;
SharedReg203_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_3_cast <= SharedReg203_out;
SharedReg43_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_4_cast <= SharedReg43_out;
   MUX_Product321_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg175_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg203_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg43_out_to_MUX_Product321_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product321_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product321_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Subtract22_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Subtract22_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Subtract22_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract22_impl_out,
                 X => Delay1No174_out_to_Subtract22_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Subtract22_impl_parent_implementedSystem_port_1_cast);

SharedReg134_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_1_cast <= SharedReg134_out;
SharedReg62_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg112_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_3_cast <= SharedReg112_out;
SharedReg136_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_4_cast <= SharedReg136_out;
   MUX_Subtract22_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg134_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg112_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg136_out_to_MUX_Subtract22_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract22_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_impl_0_out,
                 Y => Delay1No174_out);

SharedReg135_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_1_cast <= SharedReg135_out;
SharedReg94_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_2_cast <= SharedReg94_out;
SharedReg117_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_3_cast <= SharedReg117_out;
Delay2No68_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_4_cast <= Delay2No68_out;
   MUX_Subtract22_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg135_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg94_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg117_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay2No68_out_to_MUX_Subtract22_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract22_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract22_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product223_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product223_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product223_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product223_impl_out,
                 X => Delay1No176_out_to_Product223_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product223_impl_parent_implementedSystem_port_1_cast);

SharedReg225_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_1_cast <= SharedReg225_out;
SharedReg210_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_2_cast <= SharedReg210_out;
Delay22No_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_3_cast <= Delay22No_out;
SharedReg243_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
   MUX_Product223_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg225_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg210_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay22No_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Product223_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product223_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product223_impl_0_out,
                 Y => Delay1No176_out);

SharedReg150_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_1_cast <= SharedReg150_out;
SharedReg146_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
Delay3No8_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_3_cast <= Delay3No8_out;
SharedReg34_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_4_cast <= SharedReg34_out;
   MUX_Product223_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg150_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay3No8_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg34_out_to_MUX_Product223_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product223_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product223_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Subtract24_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Subtract24_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Subtract24_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract24_impl_out,
                 X => Delay1No178_out_to_Subtract24_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Subtract24_impl_parent_implementedSystem_port_1_cast);

SharedReg136_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_1_cast <= SharedReg136_out;
SharedReg101_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_2_cast <= SharedReg101_out;
Delay2No53_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_3_cast <= Delay2No53_out;
SharedReg138_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_4_cast <= SharedReg138_out;
   MUX_Subtract24_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg136_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg101_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No53_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg138_out_to_MUX_Subtract24_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract24_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_impl_0_out,
                 Y => Delay1No178_out);

SharedReg137_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_1_cast <= SharedReg137_out;
SharedReg108_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_2_cast <= SharedReg108_out;
Delay2No55_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_3_cast <= Delay2No55_out;
SharedReg144_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_4_cast <= SharedReg144_out;
   MUX_Subtract24_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg137_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg108_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No55_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg144_out_to_MUX_Subtract24_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract24_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract24_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product53_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product53_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product53_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product53_impl_out,
                 X => Delay1No180_out_to_Product53_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product53_impl_parent_implementedSystem_port_1_cast);

SharedReg151_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_1_cast <= SharedReg151_out;
SharedReg210_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_2_cast <= SharedReg210_out;
SharedReg208_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_3_cast <= SharedReg208_out;
SharedReg43_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_4_cast <= SharedReg43_out;
   MUX_Product53_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg151_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg210_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg208_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg43_out_to_MUX_Product53_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product53_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product53_impl_0_out,
                 Y => Delay1No180_out);

SharedReg225_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_1_cast <= SharedReg225_out;
SharedReg147_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg51_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_3_cast <= SharedReg51_out;
SharedReg243_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_4_cast <= SharedReg243_out;
   MUX_Product53_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg225_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg51_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Product53_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product53_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product53_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product125_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product125_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product125_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product125_impl_out,
                 X => Delay1No182_out_to_Product125_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product125_impl_parent_implementedSystem_port_1_cast);

SharedReg232_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_1_cast <= SharedReg232_out;
SharedReg211_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg208_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_3_cast <= SharedReg208_out;
SharedReg246_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_4_cast <= SharedReg246_out;
   MUX_Product125_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg232_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg208_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg246_out_to_MUX_Product125_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product125_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product125_impl_0_out,
                 Y => Delay1No182_out);

SharedReg142_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg146_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
SharedReg52_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_3_cast <= SharedReg52_out;
SharedReg151_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_4_cast <= SharedReg151_out;
   MUX_Product125_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg52_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg151_out_to_MUX_Product125_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product125_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product125_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product324_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product324_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product324_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product324_impl_out,
                 X => Delay1No184_out_to_Product324_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product324_impl_parent_implementedSystem_port_1_cast);

SharedReg232_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_1_cast <= SharedReg232_out;
SharedReg147_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg52_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_3_cast <= SharedReg52_out;
SharedReg246_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_4_cast <= SharedReg246_out;
   MUX_Product324_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg232_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg52_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg246_out_to_MUX_Product324_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product324_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_impl_0_out,
                 Y => Delay1No184_out);

SharedReg145_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg211_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_2_cast <= SharedReg211_out;
SharedReg209_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_3_cast <= SharedReg209_out;
SharedReg152_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_4_cast <= SharedReg152_out;
   MUX_Product324_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg211_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg209_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg152_out_to_MUX_Product324_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product324_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product324_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Subtract25_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Subtract25_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Subtract25_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract25_impl_out,
                 X => Delay1No186_out_to_Subtract25_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Subtract25_impl_parent_implementedSystem_port_1_cast);

SharedReg55_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_1_cast <= SharedReg55_out;
SharedReg95_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg121_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_3_cast <= SharedReg121_out;
SharedReg101_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
   MUX_Subtract25_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg55_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg121_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Subtract25_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract25_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract25_impl_0_out,
                 Y => Delay1No186_out);

SharedReg96_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_1_cast <= SharedReg96_out;
SharedReg102_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_2_cast <= SharedReg102_out;
SharedReg123_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg140_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_4_cast <= SharedReg140_out;
   MUX_Subtract25_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg96_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg102_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg123_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg140_out_to_MUX_Subtract25_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract25_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract25_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Add67_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Add67_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Add67_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add67_impl_out,
                 X => Delay1No188_out_to_Add67_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Add67_impl_parent_implementedSystem_port_1_cast);

SharedReg121_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_1_cast <= SharedReg121_out;
SharedReg138_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_2_cast <= SharedReg138_out;
   MUX_Add67_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg121_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg138_out_to_MUX_Add67_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add67_impl_0_LUT_out,
                 oMux => MUX_Add67_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add67_impl_0_out,
                 Y => Delay1No188_out);

SharedReg122_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_1_cast <= SharedReg122_out;
SharedReg139_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
   MUX_Add67_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg122_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Add67_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Add67_impl_1_LUT_out,
                 oMux => MUX_Add67_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add67_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Add68_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Add68_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Add68_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add68_impl_out,
                 X => Delay1No190_out_to_Add68_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Add68_impl_parent_implementedSystem_port_1_cast);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => Delay1No190_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Product55_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Product55_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Product55_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_impl_out,
                 X => Delay1No192_out_to_Product55_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Product55_impl_parent_implementedSystem_port_1_cast);

SharedReg233_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg204_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast <= SharedReg204_out;
SharedReg230_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_3_cast <= SharedReg230_out;
SharedReg247_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_4_cast <= SharedReg247_out;
   MUX_Product55_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg204_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg230_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg247_out_to_MUX_Product55_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_impl_0_out,
                 Y => Delay1No192_out);

SharedReg142_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg148_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast <= SharedReg148_out;
SharedReg53_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_3_cast <= SharedReg53_out;
SharedReg151_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_4_cast <= SharedReg151_out;
   MUX_Product55_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg148_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg53_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg151_out_to_MUX_Product55_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product55_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product127_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product127_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product127_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product127_impl_out,
                 X => Delay1No194_out_to_Product127_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product127_impl_parent_implementedSystem_port_1_cast);

SharedReg145_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg204_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_2_cast <= SharedReg204_out;
SharedReg230_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_3_cast <= SharedReg230_out;
SharedReg152_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_4_cast <= SharedReg152_out;
   MUX_Product127_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg204_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg230_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg152_out_to_MUX_Product127_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product127_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_impl_0_out,
                 Y => Delay1No194_out);

SharedReg233_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_1_cast <= SharedReg233_out;
SharedReg149_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_2_cast <= SharedReg149_out;
SharedReg55_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg247_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_4_cast <= SharedReg247_out;
   MUX_Product127_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg233_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg247_out_to_MUX_Product127_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product127_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product127_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Product226_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Product226_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Product226_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_impl_out,
                 X => Delay1No196_out_to_Product226_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Product226_impl_parent_implementedSystem_port_1_cast);

SharedReg218_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_1_cast <= SharedReg218_out;
SharedReg205_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg231_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_3_cast <= SharedReg231_out;
SharedReg244_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_4_cast <= SharedReg244_out;
   MUX_Product226_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg218_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg231_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_Product226_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product226_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_impl_0_out,
                 Y => Delay1No196_out);

SharedReg146_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_1_cast <= SharedReg146_out;
SharedReg148_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_2_cast <= SharedReg148_out;
SharedReg53_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_3_cast <= SharedReg53_out;
SharedReg154_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_4_cast <= SharedReg154_out;
   MUX_Product226_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg146_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg148_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg53_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg154_out_to_MUX_Product226_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product226_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product326_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product326_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product326_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_impl_out,
                 X => Delay1No198_out_to_Product326_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product326_impl_parent_implementedSystem_port_1_cast);

SharedReg218_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_1_cast <= SharedReg218_out;
SharedReg149_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_2_cast <= SharedReg149_out;
SharedReg55_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_3_cast <= SharedReg55_out;
SharedReg244_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_4_cast <= SharedReg244_out;
   MUX_Product326_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg218_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg149_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg55_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg244_out_to_MUX_Product326_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product326_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_impl_0_out,
                 Y => Delay1No198_out);

SharedReg147_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_1_cast <= SharedReg147_out;
SharedReg205_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg231_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_3_cast <= SharedReg231_out;
SharedReg156_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_4_cast <= SharedReg156_out;
   MUX_Product326_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg147_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg231_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg156_out_to_MUX_Product326_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Product326_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Subtract36_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Subtract36_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Subtract36_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract36_impl_out,
                 X => Delay1No200_out_to_Subtract36_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Subtract36_impl_parent_implementedSystem_port_1_cast);

SharedReg118_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_1_cast <= SharedReg118_out;
SharedReg1_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg127_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_3_cast <= SharedReg127_out;
SharedReg53_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_4_cast <= SharedReg53_out;
   MUX_Subtract36_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg118_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg127_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg53_out_to_MUX_Subtract36_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract36_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract36_impl_0_out,
                 Y => Delay1No200_out);

SharedReg72_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_1_cast <= SharedReg72_out;
SharedReg17_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg130_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_3_cast <= SharedReg130_out;
SharedReg94_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_4_cast <= SharedReg94_out;
   MUX_Subtract36_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg72_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg130_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg94_out_to_MUX_Subtract36_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract36_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract36_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Product237_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Product237_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Product237_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product237_impl_out,
                 X => Delay1No202_out_to_Product237_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Product237_impl_parent_implementedSystem_port_1_cast);

SharedReg219_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_1_cast <= SharedReg219_out;
SharedReg245_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_2_cast <= SharedReg245_out;
SharedReg250_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_3_cast <= SharedReg250_out;
   MUX_Product237_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg219_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg245_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg250_out_to_MUX_Product237_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product237_impl_0_LUT_out,
                 oMux => MUX_Product237_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product237_impl_0_out,
                 Y => Delay1No202_out);

SharedReg39_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_1_cast <= SharedReg39_out;
SharedReg146_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
SharedReg154_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_3_cast <= SharedReg154_out;
   MUX_Product237_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg39_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg154_out_to_MUX_Product237_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product237_impl_1_LUT_out,
                 oMux => MUX_Product237_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product237_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Product337_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Product337_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Product337_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product337_impl_out,
                 X => Delay1No204_out_to_Product337_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Product337_impl_parent_implementedSystem_port_1_cast);

SharedReg147_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_1_cast <= SharedReg147_out;
SharedReg156_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_2_cast <= SharedReg156_out;
SharedReg250_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_3_cast <= SharedReg250_out;
   MUX_Product337_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg147_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg156_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg250_out_to_MUX_Product337_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product337_impl_0_LUT_out,
                 oMux => MUX_Product337_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product337_impl_0_out,
                 Y => Delay1No204_out);

SharedReg56_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg219_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_2_cast <= SharedReg219_out;
SharedReg245_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_3_cast <= SharedReg245_out;
   MUX_Product337_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg219_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg245_out_to_MUX_Product337_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product337_impl_1_LUT_out,
                 oMux => MUX_Product337_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product337_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product67_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product67_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product67_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product67_impl_out,
                 X => Delay1No206_out_to_Product67_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product67_impl_parent_implementedSystem_port_1_cast);

Delay36No34_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_1_cast <= Delay36No34_out;
SharedReg248_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_2_cast <= SharedReg248_out;
SharedReg251_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_3_cast <= SharedReg251_out;
   MUX_Product67_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay36No34_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg248_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg251_out_to_MUX_Product67_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product67_impl_0_LUT_out,
                 oMux => MUX_Product67_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_impl_0_out,
                 Y => Delay1No206_out);

SharedReg44_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_1_cast <= SharedReg44_out;
SharedReg39_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
Delay2No72_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_3_cast <= Delay2No72_out;
   MUX_Product67_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg44_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No72_out_to_MUX_Product67_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product67_impl_1_LUT_out,
                 oMux => MUX_Product67_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product67_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product338_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product338_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product338_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product338_impl_out,
                 X => Delay1No208_out_to_Product338_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product338_impl_parent_implementedSystem_port_1_cast);

SharedReg46_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_1_cast <= SharedReg46_out;
SharedReg56_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_2_cast <= SharedReg56_out;
Delay2No73_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_3_cast <= Delay2No73_out;
   MUX_Product338_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg46_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg56_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No73_out_to_MUX_Product338_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product338_impl_0_LUT_out,
                 oMux => MUX_Product338_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product338_impl_0_out,
                 Y => Delay1No208_out);

Delay36No35_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_1_cast <= Delay36No35_out;
SharedReg249_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_2_cast <= SharedReg249_out;
SharedReg251_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_3_cast <= SharedReg251_out;
   MUX_Product338_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay36No35_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg249_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg251_out_to_MUX_Product338_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product338_impl_1_LUT_out,
                 oMux => MUX_Product338_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product338_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product68_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product68_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product68_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product68_impl_out,
                 X => Delay1No210_out_to_Product68_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product68_impl_parent_implementedSystem_port_1_cast);

Delay36No32_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_1_cast <= Delay36No32_out;
SharedReg252_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_2_cast <= SharedReg252_out;
Delay7No17_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_3_cast <= Delay7No17_out;
   MUX_Product68_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay36No32_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay7No17_out_to_MUX_Product68_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product68_impl_0_LUT_out,
                 oMux => MUX_Product68_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_impl_0_out,
                 Y => Delay1No210_out);

SharedReg58_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_1_cast <= SharedReg58_out;
SharedReg145_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_2_cast <= SharedReg145_out;
Delay2No74_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_3_cast <= Delay2No74_out;
   MUX_Product68_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg58_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No74_out_to_MUX_Product68_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product68_impl_1_LUT_out,
                 oMux => MUX_Product68_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product68_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product339_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product339_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product339_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product339_impl_out,
                 X => Delay1No212_out_to_Product339_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product339_impl_parent_implementedSystem_port_1_cast);

Delay2No75_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_1_cast <= Delay2No75_out;
SharedReg252_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_2_cast <= SharedReg252_out;
Delay7No18_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_3_cast <= Delay7No18_out;
   MUX_Product339_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No75_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg252_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay7No18_out_to_MUX_Product339_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product339_impl_0_LUT_out,
                 oMux => MUX_Product339_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product339_impl_0_out,
                 Y => Delay1No212_out);

SharedReg60_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg145_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_2_cast <= SharedReg145_out;
Delay36No33_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_3_cast <= Delay36No33_out;
   MUX_Product339_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg145_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay36No33_out_to_MUX_Product339_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product339_impl_1_LUT_out,
                 oMux => MUX_Product339_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product339_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product145_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product145_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product145_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product145_impl_out,
                 X => Delay1No214_out_to_Product145_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product145_impl_parent_implementedSystem_port_1_cast);

Delay8No3_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_1_cast <= Delay8No3_out;
SharedReg253_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_2_cast <= SharedReg253_out;
SharedReg256_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_3_cast <= SharedReg256_out;
   MUX_Product145_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay8No3_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg253_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg256_out_to_MUX_Product145_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product145_impl_0_LUT_out,
                 oMux => MUX_Product145_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product145_impl_0_out,
                 Y => Delay1No214_out);

Delay2No29_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_1_cast <= Delay2No29_out;
SharedReg58_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_2_cast <= SharedReg58_out;
SharedReg141_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_3_cast <= SharedReg141_out;
   MUX_Product145_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No29_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg58_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg141_out_to_MUX_Product145_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product145_impl_1_LUT_out,
                 oMux => MUX_Product145_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product145_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Product244_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Product244_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Product244_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product244_impl_out,
                 X => Delay1No216_out_to_Product244_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Product244_impl_parent_implementedSystem_port_1_cast);

SharedReg60_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
Delay8No4_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_2_cast <= Delay8No4_out;
SharedReg256_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_3_cast <= SharedReg256_out;
   MUX_Product244_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay8No4_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg256_out_to_MUX_Product244_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product244_impl_0_LUT_out,
                 oMux => MUX_Product244_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product244_impl_0_out,
                 Y => Delay1No216_out);

SharedReg45_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_1_cast <= SharedReg45_out;
SharedReg146_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_2_cast <= SharedReg146_out;
SharedReg253_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_3_cast <= SharedReg253_out;
   MUX_Product244_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg45_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg253_out_to_MUX_Product244_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Product244_impl_1_LUT_out,
                 oMux => MUX_Product244_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product244_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Subtract46_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Subtract46_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Subtract46_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract46_impl_out,
                 X => Delay1No218_out_to_Subtract46_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Subtract46_impl_parent_implementedSystem_port_1_cast);

SharedReg103_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_1_cast <= SharedReg103_out;
SharedReg2_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg132_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_3_cast <= SharedReg132_out;
SharedReg124_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_4_cast <= SharedReg124_out;
   MUX_Subtract46_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg103_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg132_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg124_out_to_MUX_Subtract46_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract46_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_impl_0_out,
                 Y => Delay1No218_out);

SharedReg51_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_1_cast <= SharedReg51_out;
SharedReg18_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg135_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_3_cast <= SharedReg135_out;
SharedReg142_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_4_cast <= SharedReg142_out;
   MUX_Subtract46_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg51_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg135_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg142_out_to_MUX_Subtract46_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract46_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract46_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Subtract47_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Subtract47_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Subtract47_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract47_impl_out,
                 X => Delay1No220_out_to_Subtract47_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Subtract47_impl_parent_implementedSystem_port_1_cast);

SharedReg120_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_1_cast <= SharedReg120_out;
SharedReg4_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg136_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_3_cast <= SharedReg136_out;
SharedReg88_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_4_cast <= SharedReg88_out;
   MUX_Subtract47_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg120_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg136_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg88_out_to_MUX_Subtract47_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract47_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_impl_0_out,
                 Y => Delay1No220_out);

SharedReg67_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_1_cast <= SharedReg67_out;
SharedReg20_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg139_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_3_cast <= SharedReg139_out;
SharedReg108_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_4_cast <= SharedReg108_out;
   MUX_Subtract47_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg67_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg139_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg108_out_to_MUX_Subtract47_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract47_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract47_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Product148_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Product148_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Product148_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product148_impl_out,
                 X => Delay1No222_out_to_Product148_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Product148_impl_parent_implementedSystem_port_1_cast);

SharedReg254_out_to_MUX_Product148_impl_0_parent_implementedSystem_port_1_cast <= SharedReg254_out;
SharedReg257_out_to_MUX_Product148_impl_0_parent_implementedSystem_port_2_cast <= SharedReg257_out;
   MUX_Product148_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg254_out_to_MUX_Product148_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product148_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product148_impl_0_LUT_out,
                 oMux => MUX_Product148_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product148_impl_0_out,
                 Y => Delay1No222_out);

SharedReg131_out_to_MUX_Product148_impl_1_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg141_out_to_MUX_Product148_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
   MUX_Product148_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product148_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Product148_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product148_impl_1_LUT_out,
                 oMux => MUX_Product148_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product148_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Product347_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Product347_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Product347_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product347_impl_out,
                 X => Delay1No224_out_to_Product347_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Product347_impl_parent_implementedSystem_port_1_cast);

SharedReg131_out_to_MUX_Product347_impl_0_parent_implementedSystem_port_1_cast <= SharedReg131_out;
SharedReg146_out_to_MUX_Product347_impl_0_parent_implementedSystem_port_2_cast <= SharedReg146_out;
   MUX_Product347_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg131_out_to_MUX_Product347_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg146_out_to_MUX_Product347_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product347_impl_0_LUT_out,
                 oMux => MUX_Product347_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product347_impl_0_out,
                 Y => Delay1No224_out);

SharedReg255_out_to_MUX_Product347_impl_1_parent_implementedSystem_port_1_cast <= SharedReg255_out;
SharedReg257_out_to_MUX_Product347_impl_1_parent_implementedSystem_port_2_cast <= SharedReg257_out;
   MUX_Product347_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg255_out_to_MUX_Product347_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product347_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Product347_impl_1_LUT_out,
                 oMux => MUX_Product347_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product347_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Subtract50_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Subtract50_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Subtract50_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract50_impl_out,
                 X => Delay1No226_out_to_Subtract50_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Subtract50_impl_parent_implementedSystem_port_1_cast);

SharedReg104_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_1_cast <= SharedReg104_out;
SharedReg5_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
Delay2No_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_3_cast <= Delay2No_out;
SharedReg51_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_4_cast <= SharedReg51_out;
   MUX_Subtract50_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg104_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg51_out_to_MUX_Subtract50_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract50_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract50_impl_0_out,
                 Y => Delay1No226_out);

SharedReg52_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_1_cast <= SharedReg52_out;
SharedReg21_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
Delay2No9_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_3_cast <= Delay2No9_out;
SharedReg55_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_4_cast <= SharedReg55_out;
   MUX_Subtract50_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg52_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay2No9_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg55_out_to_MUX_Subtract50_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract50_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract50_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Subtract111_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Subtract111_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Subtract111_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract111_impl_out,
                 X => Delay1No228_out_to_Subtract111_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Subtract111_impl_parent_implementedSystem_port_1_cast);

Delay2No36_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_1_cast <= Delay2No36_out;
SharedReg78_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_2_cast <= SharedReg78_out;
SharedReg3_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_3_cast <= SharedReg3_out;
SharedReg93_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_4_cast <= SharedReg93_out;
   MUX_Subtract111_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No36_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg78_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg3_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg93_out_to_MUX_Subtract111_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract111_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract111_impl_0_out,
                 Y => Delay1No228_out);

SharedReg86_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg93_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_2_cast <= SharedReg93_out;
SharedReg19_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg110_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_4_cast <= SharedReg110_out;
   MUX_Subtract111_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg93_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg19_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg110_out_to_MUX_Subtract111_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract111_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract111_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Subtract116_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Subtract116_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Subtract116_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract116_impl_out,
                 X => Delay1No230_out_to_Subtract116_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Subtract116_impl_parent_implementedSystem_port_1_cast);

SharedReg49_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_1_cast <= SharedReg49_out;
SharedReg60_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_2_cast <= SharedReg60_out;
SharedReg72_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_3_cast <= SharedReg72_out;
SharedReg52_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_4_cast <= SharedReg52_out;
   MUX_Subtract116_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg49_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg60_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg72_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg52_out_to_MUX_Subtract116_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract116_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract116_impl_0_out,
                 Y => Delay1No230_out);

Delay2No40_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_1_cast <= Delay2No40_out;
SharedReg61_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg78_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_3_cast <= SharedReg78_out;
SharedReg56_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_4_cast <= SharedReg56_out;
   MUX_Subtract116_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No40_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg78_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg56_out_to_MUX_Subtract116_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract116_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract116_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Subtract57_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Subtract57_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Subtract57_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract57_impl_out,
                 X => Delay1No232_out_to_Subtract57_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Subtract57_impl_parent_implementedSystem_port_1_cast);

SharedReg73_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_1_cast <= SharedReg73_out;
SharedReg110_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_2_cast <= SharedReg110_out;
SharedReg94_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_3_cast <= SharedReg94_out;
SharedReg113_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_4_cast <= SharedReg113_out;
   MUX_Subtract57_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg73_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg110_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg94_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg113_out_to_MUX_Subtract57_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract57_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_impl_0_out,
                 Y => Delay1No232_out);

SharedReg78_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_1_cast <= SharedReg78_out;
SharedReg113_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_2_cast <= SharedReg113_out;
SharedReg57_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_3_cast <= SharedReg57_out;
SharedReg69_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_4_cast <= SharedReg69_out;
   MUX_Subtract57_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg78_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg113_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg57_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg69_out_to_MUX_Subtract57_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract57_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract57_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Subtract117_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Subtract117_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Subtract117_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract117_impl_out,
                 X => Delay1No234_out_to_Subtract117_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Subtract117_impl_parent_implementedSystem_port_1_cast);

SharedReg50_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_1_cast <= SharedReg50_out;
Delay2No58_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_2_cast <= Delay2No58_out;
SharedReg67_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg58_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_4_cast <= SharedReg58_out;
   MUX_Subtract117_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg50_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay2No58_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg67_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg58_out_to_MUX_Subtract117_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract117_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_impl_0_out,
                 Y => Delay1No234_out);

SharedReg53_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_1_cast <= SharedReg53_out;
SharedReg86_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_2_cast <= SharedReg86_out;
SharedReg93_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_3_cast <= SharedReg93_out;
SharedReg59_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_4_cast <= SharedReg59_out;
   MUX_Subtract117_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg53_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg86_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg93_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg59_out_to_MUX_Subtract117_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract117_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract117_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Subtract61_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Subtract61_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Subtract61_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract61_impl_out,
                 X => Delay1No236_out_to_Subtract61_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Subtract61_impl_parent_implementedSystem_port_1_cast);

SharedReg56_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg118_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_2_cast <= SharedReg118_out;
SharedReg95_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg118_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_4_cast <= SharedReg118_out;
   MUX_Subtract61_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg118_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg118_out_to_MUX_Subtract61_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract61_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract61_impl_0_out,
                 Y => Delay1No236_out);

SharedReg58_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_1_cast <= SharedReg58_out;
SharedReg120_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_2_cast <= SharedReg120_out;
SharedReg102_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_3_cast <= SharedReg102_out;
SharedReg120_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_4_cast <= SharedReg120_out;
   MUX_Subtract61_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg58_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg120_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg102_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg120_out_to_MUX_Subtract61_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract61_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract61_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Subtract121_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Subtract121_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Subtract121_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract121_impl_out,
                 X => Delay1No238_out_to_Subtract121_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Subtract121_impl_parent_implementedSystem_port_1_cast);

SharedReg60_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_1_cast <= SharedReg60_out;
SharedReg6_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_2_cast <= SharedReg6_out;
SharedReg85_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_3_cast <= SharedReg85_out;
SharedReg60_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_4_cast <= SharedReg60_out;
   MUX_Subtract121_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg60_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg6_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg85_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg60_out_to_MUX_Subtract121_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract121_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract121_impl_0_out,
                 Y => Delay1No238_out);

SharedReg61_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg22_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_2_cast <= SharedReg22_out;
SharedReg101_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_3_cast <= SharedReg101_out;
SharedReg61_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_4_cast <= SharedReg61_out;
   MUX_Subtract121_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg22_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg101_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg61_out_to_MUX_Subtract121_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract121_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract121_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Subtract125_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Subtract125_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Subtract125_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract125_impl_out,
                 X => Delay1No240_out_to_Subtract125_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Subtract125_impl_parent_implementedSystem_port_1_cast);

SharedReg88_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_1_cast <= SharedReg88_out;
SharedReg7_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_2_cast <= SharedReg7_out;
SharedReg103_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_3_cast <= SharedReg103_out;
SharedReg67_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_4_cast <= SharedReg67_out;
   MUX_Subtract125_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg88_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg7_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg103_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg67_out_to_MUX_Subtract125_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract125_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract125_impl_0_out,
                 Y => Delay1No240_out);

SharedReg101_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_1_cast <= SharedReg101_out;
SharedReg23_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_2_cast <= SharedReg23_out;
SharedReg125_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_3_cast <= SharedReg125_out;
SharedReg131_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_4_cast <= SharedReg131_out;
   MUX_Subtract125_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg101_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg23_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg125_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg131_out_to_MUX_Subtract125_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract125_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract125_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Subtract66_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Subtract66_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Subtract66_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract66_impl_out,
                 X => Delay1No242_out_to_Subtract66_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Subtract66_impl_parent_implementedSystem_port_1_cast);

SharedReg62_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_1_cast <= SharedReg62_out;
SharedReg8_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_2_cast <= SharedReg8_out;
SharedReg88_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_3_cast <= SharedReg88_out;
SharedReg47_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_4_cast <= SharedReg47_out;
   MUX_Subtract66_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg62_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg8_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg88_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg47_out_to_MUX_Subtract66_impl_0_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract66_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract66_impl_0_out,
                 Y => Delay1No242_out);

SharedReg94_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_1_cast <= SharedReg94_out;
SharedReg24_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_2_cast <= SharedReg24_out;
SharedReg108_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_3_cast <= SharedReg108_out;
SharedReg62_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
   MUX_Subtract66_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg94_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg24_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg108_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Subtract66_impl_1_parent_implementedSystem_port_4_cast,
                 iSel => ModCount41_out,
                 oMux => MUX_Subtract66_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract66_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Subtract126_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Subtract126_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Subtract126_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract126_impl_out,
                 X => Delay1No244_out_to_Subtract126_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Subtract126_impl_parent_implementedSystem_port_1_cast);

SharedReg10_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_1_cast <= SharedReg10_out;
SharedReg104_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_2_cast <= SharedReg104_out;
SharedReg108_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_3_cast <= SharedReg108_out;
   MUX_Subtract126_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg10_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg104_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg108_out_to_MUX_Subtract126_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Subtract126_impl_0_LUT_out,
                 oMux => MUX_Subtract126_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract126_impl_0_out,
                 Y => Delay1No244_out);

SharedReg26_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_1_cast <= SharedReg26_out;
SharedReg126_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_2_cast <= SharedReg126_out;
SharedReg110_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_3_cast <= SharedReg110_out;
   MUX_Subtract126_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg26_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg110_out_to_MUX_Subtract126_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Subtract126_impl_1_LUT_out,
                 oMux => MUX_Subtract126_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract126_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Subtract135_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Subtract135_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Subtract135_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract135_impl_out,
                 X => Delay1No246_out_to_Subtract135_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Subtract135_impl_parent_implementedSystem_port_1_cast);

Delay2No3_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_1_cast <= Delay2No3_out;
SharedReg12_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_2_cast <= SharedReg12_out;
SharedReg95_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
   MUX_Subtract135_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No3_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg12_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg95_out_to_MUX_Subtract135_impl_0_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Subtract135_impl_0_LUT_out,
                 oMux => MUX_Subtract135_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract135_impl_0_out,
                 Y => Delay1No246_out);

Delay2No12_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_1_cast <= Delay2No12_out;
SharedReg28_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_2_cast <= SharedReg28_out;
SharedReg102_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_3_cast <= SharedReg102_out;
   MUX_Subtract135_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_3_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No12_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg28_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg102_out_to_MUX_Subtract135_impl_1_parent_implementedSystem_port_3_cast,
                 iSel => MUX_Subtract135_impl_1_LUT_out,
                 oMux => MUX_Subtract135_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract135_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Subtract137_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Subtract137_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Subtract137_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract137_impl_out,
                 X => Delay1No248_out_to_Subtract137_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Subtract137_impl_parent_implementedSystem_port_1_cast);

SharedReg11_out_to_MUX_Subtract137_impl_0_parent_implementedSystem_port_1_cast <= SharedReg11_out;
SharedReg13_out_to_MUX_Subtract137_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
   MUX_Subtract137_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg11_out_to_MUX_Subtract137_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract137_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract137_impl_0_LUT_out,
                 oMux => MUX_Subtract137_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract137_impl_0_out,
                 Y => Delay1No248_out);

SharedReg27_out_to_MUX_Subtract137_impl_1_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg29_out_to_MUX_Subtract137_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
   MUX_Subtract137_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Subtract137_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract137_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract137_impl_1_LUT_out,
                 oMux => MUX_Subtract137_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract137_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Subtract79_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Subtract79_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Subtract79_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract79_impl_out,
                 X => Delay1No250_out_to_Subtract79_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Subtract79_impl_parent_implementedSystem_port_1_cast);

Delay2No7_out_to_MUX_Subtract79_impl_0_parent_implementedSystem_port_1_cast <= Delay2No7_out;
SharedReg72_out_to_MUX_Subtract79_impl_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
   MUX_Subtract79_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No7_out_to_MUX_Subtract79_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Subtract79_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract79_impl_0_LUT_out,
                 oMux => MUX_Subtract79_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract79_impl_0_out,
                 Y => Delay1No250_out);

Delay2No16_out_to_MUX_Subtract79_impl_1_parent_implementedSystem_port_1_cast <= Delay2No16_out;
SharedReg114_out_to_MUX_Subtract79_impl_1_parent_implementedSystem_port_2_cast <= SharedReg114_out;
   MUX_Subtract79_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No16_out_to_MUX_Subtract79_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg114_out_to_MUX_Subtract79_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract79_impl_1_LUT_out,
                 oMux => MUX_Subtract79_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract79_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Subtract139_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Subtract139_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Subtract139_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract139_impl_out,
                 X => Delay1No252_out_to_Subtract139_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Subtract139_impl_parent_implementedSystem_port_1_cast);

Delay2No8_out_to_MUX_Subtract139_impl_0_parent_implementedSystem_port_1_cast <= Delay2No8_out;
SharedReg55_out_to_MUX_Subtract139_impl_0_parent_implementedSystem_port_2_cast <= SharedReg55_out;
   MUX_Subtract139_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No8_out_to_MUX_Subtract139_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg55_out_to_MUX_Subtract139_impl_0_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract139_impl_0_LUT_out,
                 oMux => MUX_Subtract139_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract139_impl_0_out,
                 Y => Delay1No252_out);

Delay2No17_out_to_MUX_Subtract139_impl_1_parent_implementedSystem_port_1_cast <= Delay2No17_out;
SharedReg125_out_to_MUX_Subtract139_impl_1_parent_implementedSystem_port_2_cast <= SharedReg125_out;
   MUX_Subtract139_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay2No17_out_to_MUX_Subtract139_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg125_out_to_MUX_Subtract139_impl_1_parent_implementedSystem_port_2_cast,
                 iSel => MUX_Subtract139_impl_1_LUT_out,
                 oMux => MUX_Subtract139_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract139_impl_1_out,
                 Y => Delay1No253_out);
   Constant2_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_impl_out);
   Constant11_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_impl_out);
   Constant3_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant3_impl_out);
   Constant12_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant12_impl_out);
   Constant4_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_impl_out);
   Constant13_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_impl_out);
   Constant5_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_impl_out);
   Constant14_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_impl_out);
   Constant6_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_impl_out);
   Constant15_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_impl_out);
   Constant7_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_impl_out);
   Constant16_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_impl_out);
   Constant8_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_impl_out);
   Constant17_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_impl_out);
   Constant9_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_impl_out);
   Constant18_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_impl_out);
   Constant10_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant10_impl_out);
   Constant19_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant19_impl_out);
   Constant20_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant20_impl_out);
   Constant110_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant110_impl_out);
   Constant21_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant21_impl_out);
   Constant111_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant111_impl_out);
   Constant22_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant22_impl_out);
   Constant112_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant112_impl_out);
   Constant23_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant23_impl_out);
   Constant113_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant113_impl_out);
   Constant24_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant24_impl_out);
   Constant114_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant114_impl_out);
   Constant25_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant25_impl_out);
   Constant115_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant115_impl_out);
   Constant26_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant26_impl_out);
   Constant116_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant116_impl_out);
   Constant27_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant27_impl_out);
   Constant117_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant117_impl_out);
   Constant28_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant28_impl_out);
   Constant118_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant118_impl_out);
   Constant29_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant29_impl_out);
   Constant119_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant119_impl_out);
   Constant30_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant30_impl_out);
   Constant120_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant120_impl_out);
   Constant31_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant31_impl_out);
   Constant121_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant121_impl_out);
   Constant32_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant32_impl_out);
   Constant122_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant122_impl_out);
   Constant33_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant33_impl_out);
   Constant123_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant123_impl_out);
   Constant34_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant34_impl_out);
   Constant124_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant124_impl_out);
   Constant35_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant35_impl_out);
   Constant125_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant125_impl_out);
   Constant36_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant36_impl_out);
   Constant126_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant126_impl_out);
   Constant37_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant37_impl_out);
   Constant127_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant127_impl_out);
   Constant38_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant38_impl_out);
   Constant128_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant128_impl_out);
   Constant39_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant39_impl_out);
   Constant129_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant129_impl_out);
   Constant40_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant40_impl_out);
   Constant130_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant130_impl_out);
   Constant41_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant41_impl_out);
   Constant131_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant131_impl_out);
   Constant42_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant42_impl_out);
   Constant132_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant132_impl_out);
   Constant43_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant43_impl_out);
   Constant133_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant133_impl_out);
   Constant44_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant44_impl_out);
   Constant134_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant134_impl_out);
   Constant45_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant45_impl_out);
   Constant135_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant135_impl_out);
   Constant46_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant46_impl_out);
   Constant136_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant136_impl_out);
   Constant47_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant47_impl_out);
   Constant137_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant137_impl_out);
   Constant48_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant48_impl_out);
   Constant138_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant138_impl_out);
   Constant49_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant49_impl_out);
   Constant139_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant139_impl_out);
   Constant50_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant50_impl_out);
   Constant140_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant140_impl_out);
   Constant51_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant51_impl_out);
   Constant141_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant141_impl_out);
   Constant52_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant52_impl_out);
   Constant142_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant142_impl_out);
   Constant53_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant53_impl_out);
   Constant143_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant143_impl_out);
   Constant54_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant54_impl_out);
   Constant144_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant144_impl_out);
   Constant55_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant55_impl_out);
   Constant145_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant145_impl_out);
   Constant56_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant56_impl_out);
   Constant146_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant146_impl_out);
   Constant57_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant57_impl_out);
   Constant147_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant147_impl_out);
   Constant_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_impl_out);
   Constant1_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_impl_out);

   Delay2No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => Delay2No_out);

   Delay3No_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => Delay3No_out);

   Delay2No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => Delay2No3_out);

   Delay2No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => Delay2No4_out);

   Delay2No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => Delay2No7_out);

   Delay2No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => Delay2No8_out);

   Delay2No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => Delay2No9_out);

   Delay3No1_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => Delay3No1_out);

   Delay2No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => Delay2No12_out);

   Delay2No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => Delay2No13_out);

   Delay2No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => Delay2No16_out);

   Delay2No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => Delay2No17_out);

   Delay2No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => Delay2No24_out);

   Delay2No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => Delay2No27_out);

   Delay2No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => Delay2No29_out);

   Delay2No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => Delay2No36_out);

   Delay2No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => Delay2No39_out);

   Delay2No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => Delay2No40_out);

   Delay2No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => Delay2No43_out);

   Delay2No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => Delay2No44_out);

   Delay3No2_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => Delay3No2_out);

   Delay2No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay2No48_out);

   Delay2No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => Delay2No49_out);

   Delay2No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => Delay2No50_out);

   Delay2No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => Delay2No51_out);

   Delay3No3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => Delay3No3_out);

   Delay2No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => Delay2No52_out);

   Delay2No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => Delay2No53_out);

   Delay2No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => Delay2No54_out);

   Delay2No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => Delay2No55_out);

   Delay2No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => Delay2No56_out);

   Delay2No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => Delay2No57_out);

   Delay2No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => Delay2No58_out);

   Delay2No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => Delay2No60_out);

   Delay2No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => Delay2No63_out);

   Delay2No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => Delay2No66_out);

   Delay2No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => Delay2No67_out);

   Delay2No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => Delay2No68_out);

   Delay3No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => Delay3No8_out);

   Delay2No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => Delay2No72_out);

   Delay2No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => Delay2No73_out);

   Delay2No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => Delay2No74_out);

   Delay2No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => Delay2No75_out);

   Delay2No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => Delay2No76_out);

   Delay3No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => Delay3No9_out);

   Delay8No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay8No2_out);

   Delay7No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => Delay7No1_out);

   Delay7No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => Delay7No2_out);

   Delay7No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => Delay7No3_out);

   Delay22No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => Delay22No_out);

   Delay22No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => Delay22No1_out);

   Delay21No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => Delay21No14_out);

   Delay21No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => Delay21No15_out);

   Delay22No6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => Delay22No6_out);

   Delay22No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => Delay22No9_out);

   Delay21No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => Delay21No31_out);

   Delay22No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => Delay22No10_out);

   Delay7No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => Delay7No14_out);

   Delay36No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => Delay36No32_out);

   Delay36No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => Delay36No33_out);

   Delay36No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => Delay36No34_out);

   Delay36No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => Delay36No35_out);

   Delay8No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => Delay8No3_out);

   Delay8No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay8No4_out);

   Delay7No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => Delay7No17_out);

   Delay7No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => Delay7No18_out);

   MUX_Add57_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add57_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add57_impl_0_LUT_out);

   MUX_Add57_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add57_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add57_impl_1_LUT_out);

   MUX_Add58_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add58_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add58_impl_0_LUT_out);

   MUX_Add58_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add58_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add58_impl_1_LUT_out);

   MUX_Add59_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add59_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add59_impl_0_LUT_out);

   MUX_Add59_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add59_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add59_impl_1_LUT_out);

   MUX_Add67_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add67_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add67_impl_0_LUT_out);

   MUX_Add67_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add67_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Add67_impl_1_LUT_out);

   MUX_Product237_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product237_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product237_impl_0_LUT_out);

   MUX_Product237_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product237_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product237_impl_1_LUT_out);

   MUX_Product337_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product337_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product337_impl_0_LUT_out);

   MUX_Product337_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product337_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product337_impl_1_LUT_out);

   MUX_Product67_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product67_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product67_impl_0_LUT_out);

   MUX_Product67_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product67_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product67_impl_1_LUT_out);

   MUX_Product338_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product338_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product338_impl_0_LUT_out);

   MUX_Product338_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product338_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product338_impl_1_LUT_out);

   MUX_Product68_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product68_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product68_impl_0_LUT_out);

   MUX_Product68_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product68_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product68_impl_1_LUT_out);

   MUX_Product339_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product339_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product339_impl_0_LUT_out);

   MUX_Product339_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product339_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product339_impl_1_LUT_out);

   MUX_Product145_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product145_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product145_impl_0_LUT_out);

   MUX_Product145_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product145_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product145_impl_1_LUT_out);

   MUX_Product244_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product244_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product244_impl_0_LUT_out);

   MUX_Product244_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product244_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product244_impl_1_LUT_out);

   MUX_Product148_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product148_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product148_impl_0_LUT_out);

   MUX_Product148_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product148_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product148_impl_1_LUT_out);

   MUX_Product347_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product347_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product347_impl_0_LUT_out);

   MUX_Product347_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product347_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Product347_impl_1_LUT_out);

   MUX_Subtract126_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract126_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract126_impl_0_LUT_out);

   MUX_Subtract126_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract126_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract126_impl_1_LUT_out);

   MUX_Subtract135_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract135_impl_0_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract135_impl_0_LUT_out);

   MUX_Subtract135_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract135_impl_1_LUT_wIn_2_wOut_2_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract135_impl_1_LUT_out);

   MUX_Subtract137_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract137_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract137_impl_0_LUT_out);

   MUX_Subtract137_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract137_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract137_impl_1_LUT_out);

   MUX_Subtract79_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract79_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract79_impl_0_LUT_out);

   MUX_Subtract79_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract79_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract79_impl_1_LUT_out);

   MUX_Subtract139_impl_0_LUT_instance: GenericLut_LUTData_MUX_Subtract139_impl_0_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract139_impl_0_LUT_out);

   MUX_Subtract139_impl_1_LUT_instance: GenericLut_LUTData_MUX_Subtract139_impl_1_LUT_wIn_2_wOut_1_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount41_out,
                 Output => MUX_Subtract139_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_impl_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add4_impl_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add6_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add15_impl_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add7_impl_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add16_impl_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_impl_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_impl_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add22_impl_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add112_impl_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add121_impl_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add33_impl_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add34_impl_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add124_impl_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add37_impl_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add127_impl_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add129_impl_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_impl_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add130_impl_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add42_impl_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add1_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_impl_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_impl_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_impl_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_impl_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_impl_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_impl_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract3_impl_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_impl_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product13_impl_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_impl_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_impl_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_impl_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product7_impl_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product8_impl_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_impl_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product17_impl_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product27_impl_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_impl_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract8_impl_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product20_impl_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract10_impl_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product30_impl_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_impl_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_impl_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_impl_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract11_impl_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add53_impl_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add54_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product42_impl_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product114_impl_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_impl_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product313_impl_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract14_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add57_impl_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add58_impl_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add59_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product118_impl_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product217_impl_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product317_impl_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract19_impl_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product219_impl_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_impl_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product49_impl_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product220_impl_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract21_impl_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product122_impl_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product221_impl_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product321_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract22_impl_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product223_impl_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract24_impl_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product53_impl_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product125_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product324_impl_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract25_impl_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add67_impl_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add68_impl_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product127_impl_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_impl_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_impl_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract36_impl_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product237_impl_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product337_impl_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product67_impl_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product338_impl_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product68_impl_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product339_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product145_impl_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product244_impl_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract46_impl_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract47_impl_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product148_impl_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product347_impl_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract50_impl_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract111_impl_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract116_impl_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract57_impl_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract117_impl_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract61_impl_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract121_impl_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract125_impl_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract66_impl_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract126_impl_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract135_impl_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract137_impl_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract79_impl_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract139_impl_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_impl_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_impl_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant3_impl_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant12_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_impl_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_impl_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_impl_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_impl_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_impl_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_impl_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_impl_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_impl_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_impl_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_impl_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_impl_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_impl_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant10_impl_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant19_impl_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant20_impl_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant110_impl_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant21_impl_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant111_impl_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant22_impl_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant112_impl_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant23_impl_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant113_impl_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant24_impl_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant114_impl_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant25_impl_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant115_impl_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant26_impl_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant116_impl_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant27_impl_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant117_impl_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant28_impl_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant118_impl_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant29_impl_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant119_impl_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant30_impl_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant120_impl_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant31_impl_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant121_impl_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant32_impl_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant122_impl_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant33_impl_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant123_impl_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant34_impl_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant124_impl_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant35_impl_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant125_impl_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant36_impl_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant126_impl_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant37_impl_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant127_impl_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant38_impl_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant128_impl_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant39_impl_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant129_impl_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant40_impl_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant130_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant41_impl_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant131_impl_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant42_impl_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant132_impl_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant43_impl_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant133_impl_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant44_impl_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant134_impl_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant45_impl_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant135_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant46_impl_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant136_impl_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant47_impl_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant137_impl_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant48_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant138_impl_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant49_impl_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant139_impl_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant50_impl_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant140_impl_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant51_impl_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant141_impl_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant52_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant142_impl_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant53_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant143_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant54_impl_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant144_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant55_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant145_impl_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant56_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant146_impl_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant57_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant147_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_impl_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_impl_out,
                 Y => SharedReg257_out);
end architecture;

